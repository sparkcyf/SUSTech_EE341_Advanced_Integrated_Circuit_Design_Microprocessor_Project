module Mux8( // @[:@3.2]
  input clock, // @[:@4.4]
  input reset, // @[:@5.4]
  input [31:0] io_int_in_0_0, // @[:@6.4]
  input [31:0] io_int_in_0_1, // @[:@6.4]
  input [31:0] io_int_in_0_2, // @[:@6.4]
  input [31:0] io_int_in_0_3, // @[:@6.4]
  input [31:0] io_int_in_0_4, // @[:@6.4]
  input [31:0] io_int_in_0_5, // @[:@6.4]
  input [31:0] io_int_in_0_6, // @[:@6.4]
  input [31:0] io_int_in_0_7, // @[:@6.4]
  input [31:0] io_int_in_1_0, // @[:@6.4]
  input [31:0] io_int_in_1_1, // @[:@6.4]
  input [31:0] io_int_in_1_2, // @[:@6.4]
  input [31:0] io_int_in_1_3, // @[:@6.4]
  input [31:0] io_int_in_1_4, // @[:@6.4]
  input [31:0] io_int_in_1_5, // @[:@6.4]
  input [31:0] io_int_in_1_6, // @[:@6.4]
  input [31:0] io_int_in_1_7, // @[:@6.4]
  input [31:0] io_int_in_2_0, // @[:@6.4]
  input [31:0] io_int_in_2_1, // @[:@6.4]
  input [31:0] io_int_in_2_2, // @[:@6.4]
  input [31:0] io_int_in_2_3, // @[:@6.4]
  input [31:0] io_int_in_2_4, // @[:@6.4]
  input [31:0] io_int_in_2_5, // @[:@6.4]
  input [31:0] io_int_in_2_6, // @[:@6.4]
  input [31:0] io_int_in_2_7, // @[:@6.4]
  input [31:0] io_int_in_3_0, // @[:@6.4]
  input [31:0] io_int_in_3_1, // @[:@6.4]
  input [31:0] io_int_in_3_2, // @[:@6.4]
  input [31:0] io_int_in_3_3, // @[:@6.4]
  input [31:0] io_int_in_3_4, // @[:@6.4]
  input [31:0] io_int_in_3_5, // @[:@6.4]
  input [31:0] io_int_in_3_6, // @[:@6.4]
  input [31:0] io_int_in_3_7, // @[:@6.4]
  input [31:0] io_int_in_4_0, // @[:@6.4]
  input [31:0] io_int_in_4_1, // @[:@6.4]
  input [31:0] io_int_in_4_2, // @[:@6.4]
  input [31:0] io_int_in_4_3, // @[:@6.4]
  input [31:0] io_int_in_4_4, // @[:@6.4]
  input [31:0] io_int_in_4_5, // @[:@6.4]
  input [31:0] io_int_in_4_6, // @[:@6.4]
  input [31:0] io_int_in_4_7, // @[:@6.4]
  input [31:0] io_int_in_5_0, // @[:@6.4]
  input [31:0] io_int_in_5_1, // @[:@6.4]
  input [31:0] io_int_in_5_2, // @[:@6.4]
  input [31:0] io_int_in_5_3, // @[:@6.4]
  input [31:0] io_int_in_5_4, // @[:@6.4]
  input [31:0] io_int_in_5_5, // @[:@6.4]
  input [31:0] io_int_in_5_6, // @[:@6.4]
  input [31:0] io_int_in_5_7, // @[:@6.4]
  input [31:0] io_int_in_6_0, // @[:@6.4]
  input [31:0] io_int_in_6_1, // @[:@6.4]
  input [31:0] io_int_in_6_2, // @[:@6.4]
  input [31:0] io_int_in_6_3, // @[:@6.4]
  input [31:0] io_int_in_6_4, // @[:@6.4]
  input [31:0] io_int_in_6_5, // @[:@6.4]
  input [31:0] io_int_in_6_6, // @[:@6.4]
  input [31:0] io_int_in_6_7, // @[:@6.4]
  input [31:0] io_int_in_7_0, // @[:@6.4]
  input [31:0] io_int_in_7_1, // @[:@6.4]
  input [31:0] io_int_in_7_2, // @[:@6.4]
  input [31:0] io_int_in_7_3, // @[:@6.4]
  input [31:0] io_int_in_7_4, // @[:@6.4]
  input [31:0] io_int_in_7_5, // @[:@6.4]
  input [31:0] io_int_in_7_6, // @[:@6.4]
  input [31:0] io_int_in_7_7, // @[:@6.4]
  input io_tag_0, // @[:@6.4]
  input io_tag_1, // @[:@6.4]
  input io_tag_2, // @[:@6.4]
  input io_tag_3, // @[:@6.4]
  input io_tag_4, // @[:@6.4]
  input io_tag_5, // @[:@6.4]
  input io_tag_6, // @[:@6.4]
  input io_tag_7, // @[:@6.4]
  output [31:0] io_choice // @[:@6.4]
);
  assign io_choice = io_int_in_0_0; // @[Mux8.scala 40:13:@8.4]
endmodule
