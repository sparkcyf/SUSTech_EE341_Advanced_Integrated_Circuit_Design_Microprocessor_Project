module MUX8( // @[:@460.2]
  input         io_in_tag_0, // @[:@463.4]
  input         io_in_tag_1, // @[:@463.4]
  input         io_in_tag_2, // @[:@463.4]
  input         io_in_tag_3, // @[:@463.4]
  input         io_in_tag_4, // @[:@463.4]
  input         io_in_tag_5, // @[:@463.4]
  input         io_in_tag_6, // @[:@463.4]
  input         io_in_tag_7, // @[:@463.4]
  output [31:0] io_choice // @[:@463.4]
);
  wire [2:0] _GEN_0; // @[MUX8.scala 58:27:@494.18]
  wire [2:0] _GEN_1; // @[MUX8.scala 56:27:@490.16]
  wire [2:0] _GEN_2; // @[MUX8.scala 54:27:@486.14]
  wire [2:0] _GEN_3; // @[MUX8.scala 52:27:@482.12]
  wire [2:0] _GEN_4; // @[MUX8.scala 50:27:@478.10]
  wire [2:0] _GEN_5; // @[MUX8.scala 48:27:@474.8]
  wire [2:0] _GEN_6; // @[MUX8.scala 46:27:@470.6]
  wire [2:0] _GEN_7; // @[MUX8.scala 44:21:@466.4]
  assign _GEN_0 = io_in_tag_7 ? 3'h7 : 3'h0; // @[MUX8.scala 58:27:@494.18]
  assign _GEN_1 = io_in_tag_6 ? 3'h6 : _GEN_0; // @[MUX8.scala 56:27:@490.16]
  assign _GEN_2 = io_in_tag_5 ? 3'h5 : _GEN_1; // @[MUX8.scala 54:27:@486.14]
  assign _GEN_3 = io_in_tag_4 ? 3'h4 : _GEN_2; // @[MUX8.scala 52:27:@482.12]
  assign _GEN_4 = io_in_tag_3 ? 3'h3 : _GEN_3; // @[MUX8.scala 50:27:@478.10]
  assign _GEN_5 = io_in_tag_2 ? 3'h2 : _GEN_4; // @[MUX8.scala 48:27:@474.8]
  assign _GEN_6 = io_in_tag_1 ? 3'h1 : _GEN_5; // @[MUX8.scala 46:27:@470.6]
  assign _GEN_7 = io_in_tag_0 ? 3'h0 : _GEN_6; // @[MUX8.scala 44:21:@466.4]
  assign io_choice = {{29'd0}, _GEN_7}; // @[MUX8.scala 42:13:@465.4 MUX8.scala 45:15:@467.6 MUX8.scala 47:15:@471.8 MUX8.scala 49:15:@475.10 MUX8.scala 51:15:@479.12 MUX8.scala 53:15:@483.14 MUX8.scala 55:15:@487.16 MUX8.scala 57:15:@491.18 MUX8.scala 59:15:@495.20 MUX8.scala 61:15:@498.20]
endmodule
module S8DP1( // @[:@501.2]
  input         clock, // @[:@502.4]
  input         reset, // @[:@503.4]
  input  [31:0] io_in_A_0, // @[:@504.4]
  input  [31:0] io_in_A_1, // @[:@504.4]
  input  [31:0] io_in_A_2, // @[:@504.4]
  input  [31:0] io_in_A_3, // @[:@504.4]
  input  [31:0] io_in_A_4, // @[:@504.4]
  input  [31:0] io_in_A_5, // @[:@504.4]
  input  [31:0] io_in_A_6, // @[:@504.4]
  input  [31:0] io_in_A_7, // @[:@504.4]
  input  [31:0] io_in_B_0, // @[:@504.4]
  input  [31:0] io_in_B_1, // @[:@504.4]
  input  [31:0] io_in_B_2, // @[:@504.4]
  input  [31:0] io_in_B_3, // @[:@504.4]
  input  [31:0] io_in_B_4, // @[:@504.4]
  input  [31:0] io_in_B_5, // @[:@504.4]
  input  [31:0] io_in_B_6, // @[:@504.4]
  input  [31:0] io_in_B_7, // @[:@504.4]
  input         io_in_tag_0, // @[:@504.4]
  input         io_in_tag_1, // @[:@504.4]
  input         io_in_tag_2, // @[:@504.4]
  input         io_in_tag_3, // @[:@504.4]
  input         io_in_tag_4, // @[:@504.4]
  input         io_in_tag_5, // @[:@504.4]
  input         io_in_tag_6, // @[:@504.4]
  input         io_in_tag_7, // @[:@504.4]
  output [31:0] io_result, // @[:@504.4]
  input         io_in_calculate, // @[:@504.4]
  output        io_out_calculate // @[:@504.4]
);
  wire  mux_io_in_tag_0; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_1; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_2; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_3; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_4; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_5; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_6; // @[S8DP1.scala 49:19:@530.4]
  wire  mux_io_in_tag_7; // @[S8DP1.scala 49:19:@530.4]
  wire [31:0] mux_io_choice; // @[S8DP1.scala 49:19:@530.4]
  reg  tag_0; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_0;
  reg  tag_1; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_1;
  reg  tag_2; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_2;
  reg  tag_3; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_3;
  reg  tag_4; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_4;
  reg  tag_5; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_5;
  reg  tag_6; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_6;
  reg  tag_7; // @[S8DP1.scala 42:20:@515.4]
  reg [31:0] _RAND_7;
  reg [31:0] acc; // @[S8DP1.scala 44:20:@526.4]
  reg [31:0] _RAND_8;
  reg  cal; // @[S8DP1.scala 46:20:@528.4]
  reg [31:0] _RAND_9;
  reg [1:0] stateReg; // @[S8DP1.scala 54:25:@541.4]
  reg [31:0] _RAND_10;
  reg [31:0] acc_temp; // @[S8DP1.scala 56:25:@542.4]
  reg [31:0] _RAND_11;
  wire  _T_236; // @[Conditional.scala 37:30:@543.4]
  wire [2:0] _T_238; // @[:@545.6]
  wire [31:0] _GEN_1; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_2; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_3; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_4; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_5; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_6; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_7; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_9; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_10; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_11; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_12; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_13; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_14; // @[S8DP1.scala 60:48:@547.6]
  wire [31:0] _GEN_15; // @[S8DP1.scala 60:48:@547.6]
  wire [63:0] _T_241; // @[S8DP1.scala 60:48:@547.6]
  wire [63:0] _GEN_71; // @[S8DP1.scala 60:23:@548.6]
  wire [64:0] _T_242; // @[S8DP1.scala 60:23:@548.6]
  wire [63:0] _T_243; // @[S8DP1.scala 60:23:@549.6]
  wire [63:0] _T_244; // @[S8DP1.scala 60:23:@550.6]
  wire  _T_245; // @[Conditional.scala 37:30:@555.6]
  wire  _GEN_16; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_17; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_18; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_19; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_20; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_21; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_22; // @[S8DP1.scala 65:26:@559.8]
  wire  _GEN_23; // @[S8DP1.scala 65:26:@559.8]
  wire  _T_251; // @[Conditional.scala 37:30:@563.8]
  wire  _T_253; // @[S8DP1.scala 69:15:@565.10]
  wire  _T_255; // @[S8DP1.scala 69:26:@566.10]
  wire  _T_256; // @[S8DP1.scala 69:23:@567.10]
  wire  _T_258; // @[S8DP1.scala 69:39:@568.10]
  wire  _T_260; // @[S8DP1.scala 69:50:@569.10]
  wire  _T_261; // @[S8DP1.scala 69:47:@570.10]
  wire  _T_262; // @[S8DP1.scala 69:35:@571.10]
  wire  _T_264; // @[S8DP1.scala 70:11:@572.10]
  wire  _T_266; // @[S8DP1.scala 70:22:@573.10]
  wire  _T_267; // @[S8DP1.scala 70:19:@574.10]
  wire  _T_269; // @[S8DP1.scala 70:35:@575.10]
  wire  _T_271; // @[S8DP1.scala 70:46:@576.10]
  wire  _T_272; // @[S8DP1.scala 70:43:@577.10]
  wire  _T_273; // @[S8DP1.scala 70:31:@578.10]
  wire  _T_274; // @[S8DP1.scala 69:60:@579.10]
  wire [1:0] _GEN_24; // @[S8DP1.scala 70:57:@580.10]
  wire  _GEN_25; // @[S8DP1.scala 70:57:@580.10]
  wire  _T_276; // @[Conditional.scala 37:30:@589.10]
  reg  _T_278; // @[S8DP1.scala 81:40:@599.12]
  reg [31:0] _RAND_12;
  wire  _T_280; // @[S8DP1.scala 81:32:@601.12]
  wire  _T_281; // @[S8DP1.scala 81:30:@602.12]
  wire  _T_282; // @[S8DP1.scala 81:70:@603.12]
  wire  _T_283; // @[S8DP1.scala 81:80:@604.12]
  wire  _T_284; // @[S8DP1.scala 81:90:@605.12]
  wire  _T_285; // @[S8DP1.scala 81:100:@606.12]
  wire  _T_286; // @[S8DP1.scala 82:16:@607.12]
  wire  _T_287; // @[S8DP1.scala 82:26:@608.12]
  wire  _T_288; // @[S8DP1.scala 82:36:@609.12]
  wire  _T_289; // @[S8DP1.scala 81:59:@610.12]
  wire [1:0] _GEN_26; // @[S8DP1.scala 83:7:@611.12]
  wire  _GEN_27; // @[S8DP1.scala 83:7:@611.12]
  wire  _GEN_28; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_29; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_30; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_31; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_32; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_33; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_34; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_35; // @[Conditional.scala 39:67:@590.10]
  wire [1:0] _GEN_36; // @[Conditional.scala 39:67:@590.10]
  wire  _GEN_37; // @[Conditional.scala 39:67:@590.10]
  wire [1:0] _GEN_38; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_39; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_40; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_41; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_42; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_43; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_44; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_45; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_46; // @[Conditional.scala 39:67:@564.8]
  wire  _GEN_47; // @[Conditional.scala 39:67:@564.8]
  wire [31:0] _GEN_48; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_49; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_50; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_51; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_52; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_53; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_54; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_55; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_56; // @[Conditional.scala 39:67:@556.6]
  wire [1:0] _GEN_57; // @[Conditional.scala 39:67:@556.6]
  wire  _GEN_58; // @[Conditional.scala 39:67:@556.6]
  wire [63:0] _GEN_59; // @[Conditional.scala 40:58:@544.4]
  wire [1:0] _GEN_60; // @[Conditional.scala 40:58:@544.4]
  wire [31:0] _GEN_61; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_62; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_63; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_64; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_65; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_66; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_67; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_68; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_69; // @[Conditional.scala 40:58:@544.4]
  wire  _GEN_70; // @[Conditional.scala 40:58:@544.4]
  wire [31:0] _GEN_72; // @[S8DP1.scala 60:16:@551.6]
  MUX8 mux ( // @[S8DP1.scala 49:19:@530.4]
    .io_in_tag_0(mux_io_in_tag_0),
    .io_in_tag_1(mux_io_in_tag_1),
    .io_in_tag_2(mux_io_in_tag_2),
    .io_in_tag_3(mux_io_in_tag_3),
    .io_in_tag_4(mux_io_in_tag_4),
    .io_in_tag_5(mux_io_in_tag_5),
    .io_in_tag_6(mux_io_in_tag_6),
    .io_in_tag_7(mux_io_in_tag_7),
    .io_choice(mux_io_choice)
  );
  assign _T_236 = 2'h0 == stateReg; // @[Conditional.scala 37:30:@543.4]
  assign _T_238 = mux_io_choice[2:0]; // @[:@545.6]
  assign _GEN_1 = 3'h1 == _T_238 ? $signed(io_in_A_1) : $signed(io_in_A_0); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_2 = 3'h2 == _T_238 ? $signed(io_in_A_2) : $signed(_GEN_1); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_3 = 3'h3 == _T_238 ? $signed(io_in_A_3) : $signed(_GEN_2); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_4 = 3'h4 == _T_238 ? $signed(io_in_A_4) : $signed(_GEN_3); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_5 = 3'h5 == _T_238 ? $signed(io_in_A_5) : $signed(_GEN_4); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_6 = 3'h6 == _T_238 ? $signed(io_in_A_6) : $signed(_GEN_5); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_7 = 3'h7 == _T_238 ? $signed(io_in_A_7) : $signed(_GEN_6); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_9 = 3'h1 == _T_238 ? $signed(io_in_B_1) : $signed(io_in_B_0); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_10 = 3'h2 == _T_238 ? $signed(io_in_B_2) : $signed(_GEN_9); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_11 = 3'h3 == _T_238 ? $signed(io_in_B_3) : $signed(_GEN_10); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_12 = 3'h4 == _T_238 ? $signed(io_in_B_4) : $signed(_GEN_11); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_13 = 3'h5 == _T_238 ? $signed(io_in_B_5) : $signed(_GEN_12); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_14 = 3'h6 == _T_238 ? $signed(io_in_B_6) : $signed(_GEN_13); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_15 = 3'h7 == _T_238 ? $signed(io_in_B_7) : $signed(_GEN_14); // @[S8DP1.scala 60:48:@547.6]
  assign _T_241 = $signed(_GEN_7) * $signed(_GEN_15); // @[S8DP1.scala 60:48:@547.6]
  assign _GEN_71 = {{32{acc[31]}},acc}; // @[S8DP1.scala 60:23:@548.6]
  assign _T_242 = $signed(_GEN_71) + $signed(_T_241); // @[S8DP1.scala 60:23:@548.6]
  assign _T_243 = _T_242[63:0]; // @[S8DP1.scala 60:23:@549.6]
  assign _T_244 = $signed(_T_243); // @[S8DP1.scala 60:23:@550.6]
  assign _T_245 = 2'h1 == stateReg; // @[Conditional.scala 37:30:@555.6]
  assign _GEN_16 = 3'h0 == _T_238 ? 1'h0 : tag_0; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_17 = 3'h1 == _T_238 ? 1'h0 : tag_1; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_18 = 3'h2 == _T_238 ? 1'h0 : tag_2; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_19 = 3'h3 == _T_238 ? 1'h0 : tag_3; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_20 = 3'h4 == _T_238 ? 1'h0 : tag_4; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_21 = 3'h5 == _T_238 ? 1'h0 : tag_5; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_22 = 3'h6 == _T_238 ? 1'h0 : tag_6; // @[S8DP1.scala 65:26:@559.8]
  assign _GEN_23 = 3'h7 == _T_238 ? 1'h0 : tag_7; // @[S8DP1.scala 65:26:@559.8]
  assign _T_251 = 2'h2 == stateReg; // @[Conditional.scala 37:30:@563.8]
  assign _T_253 = tag_0 == 1'h0; // @[S8DP1.scala 69:15:@565.10]
  assign _T_255 = tag_1 == 1'h0; // @[S8DP1.scala 69:26:@566.10]
  assign _T_256 = _T_253 & _T_255; // @[S8DP1.scala 69:23:@567.10]
  assign _T_258 = tag_2 == 1'h0; // @[S8DP1.scala 69:39:@568.10]
  assign _T_260 = tag_3 == 1'h0; // @[S8DP1.scala 69:50:@569.10]
  assign _T_261 = _T_258 & _T_260; // @[S8DP1.scala 69:47:@570.10]
  assign _T_262 = _T_256 & _T_261; // @[S8DP1.scala 69:35:@571.10]
  assign _T_264 = tag_4 == 1'h0; // @[S8DP1.scala 70:11:@572.10]
  assign _T_266 = tag_5 == 1'h0; // @[S8DP1.scala 70:22:@573.10]
  assign _T_267 = _T_264 & _T_266; // @[S8DP1.scala 70:19:@574.10]
  assign _T_269 = tag_6 == 1'h0; // @[S8DP1.scala 70:35:@575.10]
  assign _T_271 = tag_7 == 1'h0; // @[S8DP1.scala 70:46:@576.10]
  assign _T_272 = _T_269 & _T_271; // @[S8DP1.scala 70:43:@577.10]
  assign _T_273 = _T_267 & _T_272; // @[S8DP1.scala 70:31:@578.10]
  assign _T_274 = _T_262 & _T_273; // @[S8DP1.scala 69:60:@579.10]
  assign _GEN_24 = _T_274 ? 2'h3 : 2'h0; // @[S8DP1.scala 70:57:@580.10]
  assign _GEN_25 = _T_274 ? 1'h1 : cal; // @[S8DP1.scala 70:57:@580.10]
  assign _T_276 = 2'h3 == stateReg; // @[Conditional.scala 37:30:@589.10]
  assign _T_280 = _T_278 == 1'h0; // @[S8DP1.scala 81:32:@601.12]
  assign _T_281 = io_in_calculate & _T_280; // @[S8DP1.scala 81:30:@602.12]
  assign _T_282 = tag_0 | tag_1; // @[S8DP1.scala 81:70:@603.12]
  assign _T_283 = _T_282 | tag_2; // @[S8DP1.scala 81:80:@604.12]
  assign _T_284 = _T_283 | tag_3; // @[S8DP1.scala 81:90:@605.12]
  assign _T_285 = _T_284 | tag_4; // @[S8DP1.scala 81:100:@606.12]
  assign _T_286 = _T_285 | tag_5; // @[S8DP1.scala 82:16:@607.12]
  assign _T_287 = _T_286 | tag_6; // @[S8DP1.scala 82:26:@608.12]
  assign _T_288 = _T_287 | tag_7; // @[S8DP1.scala 82:36:@609.12]
  assign _T_289 = _T_281 & _T_288; // @[S8DP1.scala 81:59:@610.12]
  assign _GEN_26 = _T_289 ? 2'h0 : stateReg; // @[S8DP1.scala 83:7:@611.12]
  assign _GEN_27 = _T_289 ? 1'h0 : cal; // @[S8DP1.scala 83:7:@611.12]
  assign _GEN_28 = _T_276 ? io_in_tag_0 : tag_0; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_29 = _T_276 ? io_in_tag_1 : tag_1; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_30 = _T_276 ? io_in_tag_2 : tag_2; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_31 = _T_276 ? io_in_tag_3 : tag_3; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_32 = _T_276 ? io_in_tag_4 : tag_4; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_33 = _T_276 ? io_in_tag_5 : tag_5; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_34 = _T_276 ? io_in_tag_6 : tag_6; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_35 = _T_276 ? io_in_tag_7 : tag_7; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_36 = _T_276 ? _GEN_26 : stateReg; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_37 = _T_276 ? _GEN_27 : cal; // @[Conditional.scala 39:67:@590.10]
  assign _GEN_38 = _T_251 ? _GEN_24 : _GEN_36; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_39 = _T_251 ? _GEN_25 : _GEN_37; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_40 = _T_251 ? tag_0 : _GEN_28; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_41 = _T_251 ? tag_1 : _GEN_29; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_42 = _T_251 ? tag_2 : _GEN_30; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_43 = _T_251 ? tag_3 : _GEN_31; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_44 = _T_251 ? tag_4 : _GEN_32; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_45 = _T_251 ? tag_5 : _GEN_33; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_46 = _T_251 ? tag_6 : _GEN_34; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_47 = _T_251 ? tag_7 : _GEN_35; // @[Conditional.scala 39:67:@564.8]
  assign _GEN_48 = _T_245 ? $signed(acc_temp) : $signed(acc); // @[Conditional.scala 39:67:@556.6]
  assign _GEN_49 = _T_245 ? _GEN_16 : _GEN_40; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_50 = _T_245 ? _GEN_17 : _GEN_41; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_51 = _T_245 ? _GEN_18 : _GEN_42; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_52 = _T_245 ? _GEN_19 : _GEN_43; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_53 = _T_245 ? _GEN_20 : _GEN_44; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_54 = _T_245 ? _GEN_21 : _GEN_45; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_55 = _T_245 ? _GEN_22 : _GEN_46; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_56 = _T_245 ? _GEN_23 : _GEN_47; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_57 = _T_245 ? 2'h2 : _GEN_38; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_58 = _T_245 ? cal : _GEN_39; // @[Conditional.scala 39:67:@556.6]
  assign _GEN_59 = _T_236 ? $signed(_T_244) : $signed({{32{acc_temp[31]}},acc_temp}); // @[Conditional.scala 40:58:@544.4]
  assign _GEN_60 = _T_236 ? 2'h1 : _GEN_57; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_61 = _T_236 ? $signed(acc) : $signed(_GEN_48); // @[Conditional.scala 40:58:@544.4]
  assign _GEN_62 = _T_236 ? tag_0 : _GEN_49; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_63 = _T_236 ? tag_1 : _GEN_50; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_64 = _T_236 ? tag_2 : _GEN_51; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_65 = _T_236 ? tag_3 : _GEN_52; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_66 = _T_236 ? tag_4 : _GEN_53; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_67 = _T_236 ? tag_5 : _GEN_54; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_68 = _T_236 ? tag_6 : _GEN_55; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_69 = _T_236 ? tag_7 : _GEN_56; // @[Conditional.scala 40:58:@544.4]
  assign _GEN_70 = _T_236 ? cal : _GEN_58; // @[Conditional.scala 40:58:@544.4]
  assign io_result = acc; // @[S8DP1.scala 45:13:@527.4]
  assign io_out_calculate = cal; // @[S8DP1.scala 47:20:@529.4]
  assign mux_io_in_tag_0 = tag_0; // @[S8DP1.scala 50:17:@533.4]
  assign mux_io_in_tag_1 = tag_1; // @[S8DP1.scala 50:17:@534.4]
  assign mux_io_in_tag_2 = tag_2; // @[S8DP1.scala 50:17:@535.4]
  assign mux_io_in_tag_3 = tag_3; // @[S8DP1.scala 50:17:@536.4]
  assign mux_io_in_tag_4 = tag_4; // @[S8DP1.scala 50:17:@537.4]
  assign mux_io_in_tag_5 = tag_5; // @[S8DP1.scala 50:17:@538.4]
  assign mux_io_in_tag_6 = tag_6; // @[S8DP1.scala 50:17:@539.4]
  assign mux_io_in_tag_7 = tag_7; // @[S8DP1.scala 50:17:@540.4]
  assign _GEN_72 = _GEN_59[31:0]; // @[S8DP1.scala 60:16:@551.6]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  tag_0 = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  tag_1 = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  tag_2 = _RAND_2[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  tag_3 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  tag_4 = _RAND_4[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  tag_5 = _RAND_5[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  tag_6 = _RAND_6[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  tag_7 = _RAND_7[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  acc = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  cal = _RAND_9[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  stateReg = _RAND_10[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  acc_temp = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  _T_278 = _RAND_12[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      tag_0 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h0 == _T_238) begin
            tag_0 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_0 <= io_in_tag_0;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_1 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h1 == _T_238) begin
            tag_1 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_1 <= io_in_tag_1;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_2 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h2 == _T_238) begin
            tag_2 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_2 <= io_in_tag_2;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_3 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h3 == _T_238) begin
            tag_3 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_3 <= io_in_tag_3;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_4 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h4 == _T_238) begin
            tag_4 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_4 <= io_in_tag_4;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_5 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h5 == _T_238) begin
            tag_5 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_5 <= io_in_tag_5;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_6 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h6 == _T_238) begin
            tag_6 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_6 <= io_in_tag_6;
            end
          end
        end
      end
    end
    if (reset) begin
      tag_7 <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          if (3'h7 == _T_238) begin
            tag_7 <= 1'h0;
          end
        end else begin
          if (!(_T_251)) begin
            if (_T_276) begin
              tag_7 <= io_in_tag_7;
            end
          end
        end
      end
    end
    if (reset) begin
      acc <= 32'sh0;
    end else begin
      if (!(_T_236)) begin
        if (_T_245) begin
          acc <= acc_temp;
        end
      end
    end
    if (reset) begin
      cal <= 1'h0;
    end else begin
      if (!(_T_236)) begin
        if (!(_T_245)) begin
          if (_T_251) begin
            if (_T_274) begin
              cal <= 1'h1;
            end
          end else begin
            if (_T_276) begin
              if (_T_289) begin
                cal <= 1'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      stateReg <= 2'h3;
    end else begin
      if (_T_236) begin
        stateReg <= 2'h1;
      end else begin
        if (_T_245) begin
          stateReg <= 2'h2;
        end else begin
          if (_T_251) begin
            if (_T_274) begin
              stateReg <= 2'h3;
            end else begin
              stateReg <= 2'h0;
            end
          end else begin
            if (_T_276) begin
              if (_T_289) begin
                stateReg <= 2'h0;
              end
            end
          end
        end
      end
    end
    if (reset) begin
      acc_temp <= 32'sh0;
    end else begin
      acc_temp <= $signed(_GEN_72);
    end
    _T_278 <= io_in_calculate;
  end
endmodule
module TPU( // @[:@1716.2]
  input         clock, // @[:@1717.4]
  input         reset, // @[:@1718.4]
  input  [31:0] io_in_A_0_0, // @[:@1719.4]
  input  [31:0] io_in_A_0_1, // @[:@1719.4]
  input  [31:0] io_in_A_0_2, // @[:@1719.4]
  input  [31:0] io_in_A_0_3, // @[:@1719.4]
  input  [31:0] io_in_A_0_4, // @[:@1719.4]
  input  [31:0] io_in_A_0_5, // @[:@1719.4]
  input  [31:0] io_in_A_0_6, // @[:@1719.4]
  input  [31:0] io_in_A_0_7, // @[:@1719.4]
  input  [31:0] io_in_A_1_0, // @[:@1719.4]
  input  [31:0] io_in_A_1_1, // @[:@1719.4]
  input  [31:0] io_in_A_1_2, // @[:@1719.4]
  input  [31:0] io_in_A_1_3, // @[:@1719.4]
  input  [31:0] io_in_A_1_4, // @[:@1719.4]
  input  [31:0] io_in_A_1_5, // @[:@1719.4]
  input  [31:0] io_in_A_1_6, // @[:@1719.4]
  input  [31:0] io_in_A_1_7, // @[:@1719.4]
  input  [31:0] io_in_B_0_0, // @[:@1719.4]
  input  [31:0] io_in_B_0_1, // @[:@1719.4]
  input  [31:0] io_in_B_0_2, // @[:@1719.4]
  input  [31:0] io_in_B_0_3, // @[:@1719.4]
  input  [31:0] io_in_B_0_4, // @[:@1719.4]
  input  [31:0] io_in_B_0_5, // @[:@1719.4]
  input  [31:0] io_in_B_0_6, // @[:@1719.4]
  input  [31:0] io_in_B_0_7, // @[:@1719.4]
  input  [31:0] io_in_B_1_0, // @[:@1719.4]
  input  [31:0] io_in_B_1_1, // @[:@1719.4]
  input  [31:0] io_in_B_1_2, // @[:@1719.4]
  input  [31:0] io_in_B_1_3, // @[:@1719.4]
  input  [31:0] io_in_B_1_4, // @[:@1719.4]
  input  [31:0] io_in_B_1_5, // @[:@1719.4]
  input  [31:0] io_in_B_1_6, // @[:@1719.4]
  input  [31:0] io_in_B_1_7, // @[:@1719.4]
  input  [31:0] io_in_B_2_0, // @[:@1719.4]
  input  [31:0] io_in_B_2_1, // @[:@1719.4]
  input  [31:0] io_in_B_2_2, // @[:@1719.4]
  input  [31:0] io_in_B_2_3, // @[:@1719.4]
  input  [31:0] io_in_B_2_4, // @[:@1719.4]
  input  [31:0] io_in_B_2_5, // @[:@1719.4]
  input  [31:0] io_in_B_2_6, // @[:@1719.4]
  input  [31:0] io_in_B_2_7, // @[:@1719.4]
  input  [31:0] io_in_B_3_0, // @[:@1719.4]
  input  [31:0] io_in_B_3_1, // @[:@1719.4]
  input  [31:0] io_in_B_3_2, // @[:@1719.4]
  input  [31:0] io_in_B_3_3, // @[:@1719.4]
  input  [31:0] io_in_B_3_4, // @[:@1719.4]
  input  [31:0] io_in_B_3_5, // @[:@1719.4]
  input  [31:0] io_in_B_3_6, // @[:@1719.4]
  input  [31:0] io_in_B_3_7, // @[:@1719.4]
  input         io_in_tag_0_0, // @[:@1719.4]
  input         io_in_tag_0_1, // @[:@1719.4]
  input         io_in_tag_0_2, // @[:@1719.4]
  input         io_in_tag_0_3, // @[:@1719.4]
  input         io_in_tag_0_4, // @[:@1719.4]
  input         io_in_tag_0_5, // @[:@1719.4]
  input         io_in_tag_0_6, // @[:@1719.4]
  input         io_in_tag_0_7, // @[:@1719.4]
  input         io_in_tag_1_0, // @[:@1719.4]
  input         io_in_tag_1_1, // @[:@1719.4]
  input         io_in_tag_1_2, // @[:@1719.4]
  input         io_in_tag_1_3, // @[:@1719.4]
  input         io_in_tag_1_4, // @[:@1719.4]
  input         io_in_tag_1_5, // @[:@1719.4]
  input         io_in_tag_1_6, // @[:@1719.4]
  input         io_in_tag_1_7, // @[:@1719.4]
  input         io_in_tag_2_0, // @[:@1719.4]
  input         io_in_tag_2_1, // @[:@1719.4]
  input         io_in_tag_2_2, // @[:@1719.4]
  input         io_in_tag_2_3, // @[:@1719.4]
  input         io_in_tag_2_4, // @[:@1719.4]
  input         io_in_tag_2_5, // @[:@1719.4]
  input         io_in_tag_2_6, // @[:@1719.4]
  input         io_in_tag_2_7, // @[:@1719.4]
  input         io_in_tag_3_0, // @[:@1719.4]
  input         io_in_tag_3_1, // @[:@1719.4]
  input         io_in_tag_3_2, // @[:@1719.4]
  input         io_in_tag_3_3, // @[:@1719.4]
  input         io_in_tag_3_4, // @[:@1719.4]
  input         io_in_tag_3_5, // @[:@1719.4]
  input         io_in_tag_3_6, // @[:@1719.4]
  input         io_in_tag_3_7, // @[:@1719.4]
  input         io_in_cal, // @[:@1719.4]
  output [31:0] io_out_A_0_0, // @[:@1719.4]
  output [31:0] io_out_A_0_1, // @[:@1719.4]
  output [31:0] io_out_A_0_2, // @[:@1719.4]
  output [31:0] io_out_A_0_3, // @[:@1719.4]
  output [31:0] io_out_A_0_4, // @[:@1719.4]
  output [31:0] io_out_A_0_5, // @[:@1719.4]
  output [31:0] io_out_A_0_6, // @[:@1719.4]
  output [31:0] io_out_A_0_7, // @[:@1719.4]
  output [31:0] io_out_A_1_0, // @[:@1719.4]
  output [31:0] io_out_A_1_1, // @[:@1719.4]
  output [31:0] io_out_A_1_2, // @[:@1719.4]
  output [31:0] io_out_A_1_3, // @[:@1719.4]
  output [31:0] io_out_A_1_4, // @[:@1719.4]
  output [31:0] io_out_A_1_5, // @[:@1719.4]
  output [31:0] io_out_A_1_6, // @[:@1719.4]
  output [31:0] io_out_A_1_7, // @[:@1719.4]
  output [31:0] io_out_B_0_0, // @[:@1719.4]
  output [31:0] io_out_B_0_1, // @[:@1719.4]
  output [31:0] io_out_B_0_2, // @[:@1719.4]
  output [31:0] io_out_B_0_3, // @[:@1719.4]
  output [31:0] io_out_B_0_4, // @[:@1719.4]
  output [31:0] io_out_B_0_5, // @[:@1719.4]
  output [31:0] io_out_B_0_6, // @[:@1719.4]
  output [31:0] io_out_B_0_7, // @[:@1719.4]
  output [31:0] io_out_B_1_0, // @[:@1719.4]
  output [31:0] io_out_B_1_1, // @[:@1719.4]
  output [31:0] io_out_B_1_2, // @[:@1719.4]
  output [31:0] io_out_B_1_3, // @[:@1719.4]
  output [31:0] io_out_B_1_4, // @[:@1719.4]
  output [31:0] io_out_B_1_5, // @[:@1719.4]
  output [31:0] io_out_B_1_6, // @[:@1719.4]
  output [31:0] io_out_B_1_7, // @[:@1719.4]
  output [31:0] io_out_B_2_0, // @[:@1719.4]
  output [31:0] io_out_B_2_1, // @[:@1719.4]
  output [31:0] io_out_B_2_2, // @[:@1719.4]
  output [31:0] io_out_B_2_3, // @[:@1719.4]
  output [31:0] io_out_B_2_4, // @[:@1719.4]
  output [31:0] io_out_B_2_5, // @[:@1719.4]
  output [31:0] io_out_B_2_6, // @[:@1719.4]
  output [31:0] io_out_B_2_7, // @[:@1719.4]
  output [31:0] io_out_B_3_0, // @[:@1719.4]
  output [31:0] io_out_B_3_1, // @[:@1719.4]
  output [31:0] io_out_B_3_2, // @[:@1719.4]
  output [31:0] io_out_B_3_3, // @[:@1719.4]
  output [31:0] io_out_B_3_4, // @[:@1719.4]
  output [31:0] io_out_B_3_5, // @[:@1719.4]
  output [31:0] io_out_B_3_6, // @[:@1719.4]
  output [31:0] io_out_B_3_7, // @[:@1719.4]
  output        io_out_tag_0_0, // @[:@1719.4]
  output        io_out_tag_0_1, // @[:@1719.4]
  output        io_out_tag_0_2, // @[:@1719.4]
  output        io_out_tag_0_3, // @[:@1719.4]
  output        io_out_tag_0_4, // @[:@1719.4]
  output        io_out_tag_0_5, // @[:@1719.4]
  output        io_out_tag_0_6, // @[:@1719.4]
  output        io_out_tag_0_7, // @[:@1719.4]
  output        io_out_tag_1_0, // @[:@1719.4]
  output        io_out_tag_1_1, // @[:@1719.4]
  output        io_out_tag_1_2, // @[:@1719.4]
  output        io_out_tag_1_3, // @[:@1719.4]
  output        io_out_tag_1_4, // @[:@1719.4]
  output        io_out_tag_1_5, // @[:@1719.4]
  output        io_out_tag_1_6, // @[:@1719.4]
  output        io_out_tag_1_7, // @[:@1719.4]
  output        io_out_tag_2_0, // @[:@1719.4]
  output        io_out_tag_2_1, // @[:@1719.4]
  output        io_out_tag_2_2, // @[:@1719.4]
  output        io_out_tag_2_3, // @[:@1719.4]
  output        io_out_tag_2_4, // @[:@1719.4]
  output        io_out_tag_2_5, // @[:@1719.4]
  output        io_out_tag_2_6, // @[:@1719.4]
  output        io_out_tag_2_7, // @[:@1719.4]
  output        io_out_tag_3_0, // @[:@1719.4]
  output        io_out_tag_3_1, // @[:@1719.4]
  output        io_out_tag_3_2, // @[:@1719.4]
  output        io_out_tag_3_3, // @[:@1719.4]
  output        io_out_tag_3_4, // @[:@1719.4]
  output        io_out_tag_3_5, // @[:@1719.4]
  output        io_out_tag_3_6, // @[:@1719.4]
  output        io_out_tag_3_7, // @[:@1719.4]
  output [31:0] io_out_result_0_0, // @[:@1719.4]
  output [31:0] io_out_result_0_1, // @[:@1719.4]
  output [31:0] io_out_result_0_2, // @[:@1719.4]
  output [31:0] io_out_result_0_3, // @[:@1719.4]
  output [31:0] io_out_result_1_0, // @[:@1719.4]
  output [31:0] io_out_result_1_1, // @[:@1719.4]
  output [31:0] io_out_result_1_2, // @[:@1719.4]
  output [31:0] io_out_result_1_3, // @[:@1719.4]
  output        io_out_cal // @[:@1719.4]
);
  wire  S8DP1_clock; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_reset; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_0; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_1; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_2; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_3; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_4; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_5; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_6; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_A_7; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_0; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_1; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_2; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_3; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_4; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_5; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_6; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_in_B_7; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_0; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_1; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_2; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_3; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_4; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_5; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_6; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_tag_7; // @[TPU.scala 62:39:@1801.4]
  wire [31:0] S8DP1_io_result; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_in_calculate; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_io_out_calculate; // @[TPU.scala 62:39:@1801.4]
  wire  S8DP1_1_clock; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_reset; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_0; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_1; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_2; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_3; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_4; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_5; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_6; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_A_7; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_0; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_1; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_2; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_3; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_4; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_5; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_6; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_in_B_7; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_0; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_1; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_2; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_3; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_4; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_5; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_6; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_tag_7; // @[TPU.scala 62:39:@1804.4]
  wire [31:0] S8DP1_1_io_result; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_in_calculate; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_1_io_out_calculate; // @[TPU.scala 62:39:@1804.4]
  wire  S8DP1_2_clock; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_reset; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_0; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_1; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_2; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_3; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_4; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_5; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_6; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_A_7; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_0; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_1; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_2; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_3; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_4; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_5; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_6; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_in_B_7; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_0; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_1; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_2; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_3; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_4; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_5; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_6; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_tag_7; // @[TPU.scala 62:39:@1807.4]
  wire [31:0] S8DP1_2_io_result; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_in_calculate; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_2_io_out_calculate; // @[TPU.scala 62:39:@1807.4]
  wire  S8DP1_3_clock; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_reset; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_0; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_1; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_2; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_3; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_4; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_5; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_6; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_A_7; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_0; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_1; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_2; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_3; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_4; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_5; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_6; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_in_B_7; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_0; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_1; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_2; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_3; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_4; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_5; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_6; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_tag_7; // @[TPU.scala 62:39:@1810.4]
  wire [31:0] S8DP1_3_io_result; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_in_calculate; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_3_io_out_calculate; // @[TPU.scala 62:39:@1810.4]
  wire  S8DP1_4_clock; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_reset; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_0; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_1; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_2; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_3; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_4; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_5; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_6; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_A_7; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_0; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_1; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_2; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_3; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_4; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_5; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_6; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_in_B_7; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_0; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_1; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_2; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_3; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_4; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_5; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_6; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_tag_7; // @[TPU.scala 63:39:@1922.4]
  wire [31:0] S8DP1_4_io_result; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_in_calculate; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_4_io_out_calculate; // @[TPU.scala 63:39:@1922.4]
  wire  S8DP1_5_clock; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_reset; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_0; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_1; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_2; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_3; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_4; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_5; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_6; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_A_7; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_0; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_1; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_2; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_3; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_4; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_5; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_6; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_in_B_7; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_0; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_1; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_2; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_3; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_4; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_5; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_6; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_tag_7; // @[TPU.scala 63:39:@1925.4]
  wire [31:0] S8DP1_5_io_result; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_in_calculate; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_5_io_out_calculate; // @[TPU.scala 63:39:@1925.4]
  wire  S8DP1_6_clock; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_reset; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_0; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_1; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_2; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_3; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_4; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_5; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_6; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_A_7; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_0; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_1; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_2; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_3; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_4; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_5; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_6; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_in_B_7; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_0; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_1; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_2; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_3; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_4; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_5; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_6; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_tag_7; // @[TPU.scala 63:39:@1928.4]
  wire [31:0] S8DP1_6_io_result; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_in_calculate; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_6_io_out_calculate; // @[TPU.scala 63:39:@1928.4]
  wire  S8DP1_7_clock; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_reset; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_0; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_1; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_2; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_3; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_4; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_5; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_6; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_A_7; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_0; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_1; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_2; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_3; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_4; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_5; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_6; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_in_B_7; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_0; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_1; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_2; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_3; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_4; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_5; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_6; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_tag_7; // @[TPU.scala 63:39:@1931.4]
  wire [31:0] S8DP1_7_io_result; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_in_calculate; // @[TPU.scala 63:39:@1931.4]
  wire  S8DP1_7_io_out_calculate; // @[TPU.scala 63:39:@1931.4]
  reg  cal_state; // @[TPU.scala 64:26:@2043.4]
  reg [31:0] _RAND_0;
  reg  cal_control; // @[TPU.scala 65:28:@2044.4]
  reg [31:0] _RAND_1;
  wire  S8DP1_1_1_0_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1814.4]
  wire  S8DP1_1_1_1_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1841.4]
  wire  _T_3683; // @[TPU.scala 78:42:@2245.4]
  wire  S8DP1_1_1_2_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1868.4]
  wire  _T_3684; // @[TPU.scala 78:70:@2246.4]
  wire  S8DP1_1_1_3_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1895.4]
  wire  _T_3685; // @[TPU.scala 78:98:@2247.4]
  wire  S8DP1_2_1_0_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1935.4]
  wire  _T_3686; // @[TPU.scala 79:5:@2248.4]
  wire  S8DP1_2_1_1_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1962.4]
  wire  _T_3687; // @[TPU.scala 79:33:@2249.4]
  wire  S8DP1_2_1_2_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1989.4]
  wire  _T_3688; // @[TPU.scala 79:61:@2250.4]
  wire  S8DP1_2_1_3_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@2016.4]
  wire  _T_3689; // @[TPU.scala 79:89:@2251.4]
  reg [1:0] stateReg; // @[TPU.scala 90:25:@2262.4]
  reg [31:0] _RAND_2;
  wire  _T_3691; // @[Conditional.scala 37:30:@2263.4]
  reg  _T_3693; // @[TPU.scala 93:33:@2265.6]
  reg [31:0] _RAND_3;
  wire  _T_3695; // @[TPU.scala 93:25:@2267.6]
  wire  _T_3696; // @[TPU.scala 93:23:@2268.6]
  wire [1:0] _GEN_0; // @[TPU.scala 93:46:@2269.6]
  wire  _T_3697; // @[Conditional.scala 37:30:@2274.6]
  wire  _T_3698; // @[Conditional.scala 37:30:@2279.8]
  wire [1:0] _GEN_1; // @[TPU.scala 106:23:@2282.10]
  wire  _GEN_2; // @[TPU.scala 106:23:@2282.10]
  wire  _GEN_3; // @[Conditional.scala 39:67:@2280.8]
  wire [1:0] _GEN_4; // @[Conditional.scala 39:67:@2280.8]
  wire [1:0] _GEN_5; // @[Conditional.scala 39:67:@2275.6]
  wire  _GEN_6; // @[Conditional.scala 39:67:@2275.6]
  wire [1:0] _GEN_7; // @[Conditional.scala 40:58:@2264.4]
  wire  _GEN_8; // @[Conditional.scala 40:58:@2264.4]
  S8DP1 S8DP1 ( // @[TPU.scala 62:39:@1801.4]
    .clock(S8DP1_clock),
    .reset(S8DP1_reset),
    .io_in_A_0(S8DP1_io_in_A_0),
    .io_in_A_1(S8DP1_io_in_A_1),
    .io_in_A_2(S8DP1_io_in_A_2),
    .io_in_A_3(S8DP1_io_in_A_3),
    .io_in_A_4(S8DP1_io_in_A_4),
    .io_in_A_5(S8DP1_io_in_A_5),
    .io_in_A_6(S8DP1_io_in_A_6),
    .io_in_A_7(S8DP1_io_in_A_7),
    .io_in_B_0(S8DP1_io_in_B_0),
    .io_in_B_1(S8DP1_io_in_B_1),
    .io_in_B_2(S8DP1_io_in_B_2),
    .io_in_B_3(S8DP1_io_in_B_3),
    .io_in_B_4(S8DP1_io_in_B_4),
    .io_in_B_5(S8DP1_io_in_B_5),
    .io_in_B_6(S8DP1_io_in_B_6),
    .io_in_B_7(S8DP1_io_in_B_7),
    .io_in_tag_0(S8DP1_io_in_tag_0),
    .io_in_tag_1(S8DP1_io_in_tag_1),
    .io_in_tag_2(S8DP1_io_in_tag_2),
    .io_in_tag_3(S8DP1_io_in_tag_3),
    .io_in_tag_4(S8DP1_io_in_tag_4),
    .io_in_tag_5(S8DP1_io_in_tag_5),
    .io_in_tag_6(S8DP1_io_in_tag_6),
    .io_in_tag_7(S8DP1_io_in_tag_7),
    .io_result(S8DP1_io_result),
    .io_in_calculate(S8DP1_io_in_calculate),
    .io_out_calculate(S8DP1_io_out_calculate)
  );
  S8DP1 S8DP1_1 ( // @[TPU.scala 62:39:@1804.4]
    .clock(S8DP1_1_clock),
    .reset(S8DP1_1_reset),
    .io_in_A_0(S8DP1_1_io_in_A_0),
    .io_in_A_1(S8DP1_1_io_in_A_1),
    .io_in_A_2(S8DP1_1_io_in_A_2),
    .io_in_A_3(S8DP1_1_io_in_A_3),
    .io_in_A_4(S8DP1_1_io_in_A_4),
    .io_in_A_5(S8DP1_1_io_in_A_5),
    .io_in_A_6(S8DP1_1_io_in_A_6),
    .io_in_A_7(S8DP1_1_io_in_A_7),
    .io_in_B_0(S8DP1_1_io_in_B_0),
    .io_in_B_1(S8DP1_1_io_in_B_1),
    .io_in_B_2(S8DP1_1_io_in_B_2),
    .io_in_B_3(S8DP1_1_io_in_B_3),
    .io_in_B_4(S8DP1_1_io_in_B_4),
    .io_in_B_5(S8DP1_1_io_in_B_5),
    .io_in_B_6(S8DP1_1_io_in_B_6),
    .io_in_B_7(S8DP1_1_io_in_B_7),
    .io_in_tag_0(S8DP1_1_io_in_tag_0),
    .io_in_tag_1(S8DP1_1_io_in_tag_1),
    .io_in_tag_2(S8DP1_1_io_in_tag_2),
    .io_in_tag_3(S8DP1_1_io_in_tag_3),
    .io_in_tag_4(S8DP1_1_io_in_tag_4),
    .io_in_tag_5(S8DP1_1_io_in_tag_5),
    .io_in_tag_6(S8DP1_1_io_in_tag_6),
    .io_in_tag_7(S8DP1_1_io_in_tag_7),
    .io_result(S8DP1_1_io_result),
    .io_in_calculate(S8DP1_1_io_in_calculate),
    .io_out_calculate(S8DP1_1_io_out_calculate)
  );
  S8DP1 S8DP1_2 ( // @[TPU.scala 62:39:@1807.4]
    .clock(S8DP1_2_clock),
    .reset(S8DP1_2_reset),
    .io_in_A_0(S8DP1_2_io_in_A_0),
    .io_in_A_1(S8DP1_2_io_in_A_1),
    .io_in_A_2(S8DP1_2_io_in_A_2),
    .io_in_A_3(S8DP1_2_io_in_A_3),
    .io_in_A_4(S8DP1_2_io_in_A_4),
    .io_in_A_5(S8DP1_2_io_in_A_5),
    .io_in_A_6(S8DP1_2_io_in_A_6),
    .io_in_A_7(S8DP1_2_io_in_A_7),
    .io_in_B_0(S8DP1_2_io_in_B_0),
    .io_in_B_1(S8DP1_2_io_in_B_1),
    .io_in_B_2(S8DP1_2_io_in_B_2),
    .io_in_B_3(S8DP1_2_io_in_B_3),
    .io_in_B_4(S8DP1_2_io_in_B_4),
    .io_in_B_5(S8DP1_2_io_in_B_5),
    .io_in_B_6(S8DP1_2_io_in_B_6),
    .io_in_B_7(S8DP1_2_io_in_B_7),
    .io_in_tag_0(S8DP1_2_io_in_tag_0),
    .io_in_tag_1(S8DP1_2_io_in_tag_1),
    .io_in_tag_2(S8DP1_2_io_in_tag_2),
    .io_in_tag_3(S8DP1_2_io_in_tag_3),
    .io_in_tag_4(S8DP1_2_io_in_tag_4),
    .io_in_tag_5(S8DP1_2_io_in_tag_5),
    .io_in_tag_6(S8DP1_2_io_in_tag_6),
    .io_in_tag_7(S8DP1_2_io_in_tag_7),
    .io_result(S8DP1_2_io_result),
    .io_in_calculate(S8DP1_2_io_in_calculate),
    .io_out_calculate(S8DP1_2_io_out_calculate)
  );
  S8DP1 S8DP1_3 ( // @[TPU.scala 62:39:@1810.4]
    .clock(S8DP1_3_clock),
    .reset(S8DP1_3_reset),
    .io_in_A_0(S8DP1_3_io_in_A_0),
    .io_in_A_1(S8DP1_3_io_in_A_1),
    .io_in_A_2(S8DP1_3_io_in_A_2),
    .io_in_A_3(S8DP1_3_io_in_A_3),
    .io_in_A_4(S8DP1_3_io_in_A_4),
    .io_in_A_5(S8DP1_3_io_in_A_5),
    .io_in_A_6(S8DP1_3_io_in_A_6),
    .io_in_A_7(S8DP1_3_io_in_A_7),
    .io_in_B_0(S8DP1_3_io_in_B_0),
    .io_in_B_1(S8DP1_3_io_in_B_1),
    .io_in_B_2(S8DP1_3_io_in_B_2),
    .io_in_B_3(S8DP1_3_io_in_B_3),
    .io_in_B_4(S8DP1_3_io_in_B_4),
    .io_in_B_5(S8DP1_3_io_in_B_5),
    .io_in_B_6(S8DP1_3_io_in_B_6),
    .io_in_B_7(S8DP1_3_io_in_B_7),
    .io_in_tag_0(S8DP1_3_io_in_tag_0),
    .io_in_tag_1(S8DP1_3_io_in_tag_1),
    .io_in_tag_2(S8DP1_3_io_in_tag_2),
    .io_in_tag_3(S8DP1_3_io_in_tag_3),
    .io_in_tag_4(S8DP1_3_io_in_tag_4),
    .io_in_tag_5(S8DP1_3_io_in_tag_5),
    .io_in_tag_6(S8DP1_3_io_in_tag_6),
    .io_in_tag_7(S8DP1_3_io_in_tag_7),
    .io_result(S8DP1_3_io_result),
    .io_in_calculate(S8DP1_3_io_in_calculate),
    .io_out_calculate(S8DP1_3_io_out_calculate)
  );
  S8DP1 S8DP1_4 ( // @[TPU.scala 63:39:@1922.4]
    .clock(S8DP1_4_clock),
    .reset(S8DP1_4_reset),
    .io_in_A_0(S8DP1_4_io_in_A_0),
    .io_in_A_1(S8DP1_4_io_in_A_1),
    .io_in_A_2(S8DP1_4_io_in_A_2),
    .io_in_A_3(S8DP1_4_io_in_A_3),
    .io_in_A_4(S8DP1_4_io_in_A_4),
    .io_in_A_5(S8DP1_4_io_in_A_5),
    .io_in_A_6(S8DP1_4_io_in_A_6),
    .io_in_A_7(S8DP1_4_io_in_A_7),
    .io_in_B_0(S8DP1_4_io_in_B_0),
    .io_in_B_1(S8DP1_4_io_in_B_1),
    .io_in_B_2(S8DP1_4_io_in_B_2),
    .io_in_B_3(S8DP1_4_io_in_B_3),
    .io_in_B_4(S8DP1_4_io_in_B_4),
    .io_in_B_5(S8DP1_4_io_in_B_5),
    .io_in_B_6(S8DP1_4_io_in_B_6),
    .io_in_B_7(S8DP1_4_io_in_B_7),
    .io_in_tag_0(S8DP1_4_io_in_tag_0),
    .io_in_tag_1(S8DP1_4_io_in_tag_1),
    .io_in_tag_2(S8DP1_4_io_in_tag_2),
    .io_in_tag_3(S8DP1_4_io_in_tag_3),
    .io_in_tag_4(S8DP1_4_io_in_tag_4),
    .io_in_tag_5(S8DP1_4_io_in_tag_5),
    .io_in_tag_6(S8DP1_4_io_in_tag_6),
    .io_in_tag_7(S8DP1_4_io_in_tag_7),
    .io_result(S8DP1_4_io_result),
    .io_in_calculate(S8DP1_4_io_in_calculate),
    .io_out_calculate(S8DP1_4_io_out_calculate)
  );
  S8DP1 S8DP1_5 ( // @[TPU.scala 63:39:@1925.4]
    .clock(S8DP1_5_clock),
    .reset(S8DP1_5_reset),
    .io_in_A_0(S8DP1_5_io_in_A_0),
    .io_in_A_1(S8DP1_5_io_in_A_1),
    .io_in_A_2(S8DP1_5_io_in_A_2),
    .io_in_A_3(S8DP1_5_io_in_A_3),
    .io_in_A_4(S8DP1_5_io_in_A_4),
    .io_in_A_5(S8DP1_5_io_in_A_5),
    .io_in_A_6(S8DP1_5_io_in_A_6),
    .io_in_A_7(S8DP1_5_io_in_A_7),
    .io_in_B_0(S8DP1_5_io_in_B_0),
    .io_in_B_1(S8DP1_5_io_in_B_1),
    .io_in_B_2(S8DP1_5_io_in_B_2),
    .io_in_B_3(S8DP1_5_io_in_B_3),
    .io_in_B_4(S8DP1_5_io_in_B_4),
    .io_in_B_5(S8DP1_5_io_in_B_5),
    .io_in_B_6(S8DP1_5_io_in_B_6),
    .io_in_B_7(S8DP1_5_io_in_B_7),
    .io_in_tag_0(S8DP1_5_io_in_tag_0),
    .io_in_tag_1(S8DP1_5_io_in_tag_1),
    .io_in_tag_2(S8DP1_5_io_in_tag_2),
    .io_in_tag_3(S8DP1_5_io_in_tag_3),
    .io_in_tag_4(S8DP1_5_io_in_tag_4),
    .io_in_tag_5(S8DP1_5_io_in_tag_5),
    .io_in_tag_6(S8DP1_5_io_in_tag_6),
    .io_in_tag_7(S8DP1_5_io_in_tag_7),
    .io_result(S8DP1_5_io_result),
    .io_in_calculate(S8DP1_5_io_in_calculate),
    .io_out_calculate(S8DP1_5_io_out_calculate)
  );
  S8DP1 S8DP1_6 ( // @[TPU.scala 63:39:@1928.4]
    .clock(S8DP1_6_clock),
    .reset(S8DP1_6_reset),
    .io_in_A_0(S8DP1_6_io_in_A_0),
    .io_in_A_1(S8DP1_6_io_in_A_1),
    .io_in_A_2(S8DP1_6_io_in_A_2),
    .io_in_A_3(S8DP1_6_io_in_A_3),
    .io_in_A_4(S8DP1_6_io_in_A_4),
    .io_in_A_5(S8DP1_6_io_in_A_5),
    .io_in_A_6(S8DP1_6_io_in_A_6),
    .io_in_A_7(S8DP1_6_io_in_A_7),
    .io_in_B_0(S8DP1_6_io_in_B_0),
    .io_in_B_1(S8DP1_6_io_in_B_1),
    .io_in_B_2(S8DP1_6_io_in_B_2),
    .io_in_B_3(S8DP1_6_io_in_B_3),
    .io_in_B_4(S8DP1_6_io_in_B_4),
    .io_in_B_5(S8DP1_6_io_in_B_5),
    .io_in_B_6(S8DP1_6_io_in_B_6),
    .io_in_B_7(S8DP1_6_io_in_B_7),
    .io_in_tag_0(S8DP1_6_io_in_tag_0),
    .io_in_tag_1(S8DP1_6_io_in_tag_1),
    .io_in_tag_2(S8DP1_6_io_in_tag_2),
    .io_in_tag_3(S8DP1_6_io_in_tag_3),
    .io_in_tag_4(S8DP1_6_io_in_tag_4),
    .io_in_tag_5(S8DP1_6_io_in_tag_5),
    .io_in_tag_6(S8DP1_6_io_in_tag_6),
    .io_in_tag_7(S8DP1_6_io_in_tag_7),
    .io_result(S8DP1_6_io_result),
    .io_in_calculate(S8DP1_6_io_in_calculate),
    .io_out_calculate(S8DP1_6_io_out_calculate)
  );
  S8DP1 S8DP1_7 ( // @[TPU.scala 63:39:@1931.4]
    .clock(S8DP1_7_clock),
    .reset(S8DP1_7_reset),
    .io_in_A_0(S8DP1_7_io_in_A_0),
    .io_in_A_1(S8DP1_7_io_in_A_1),
    .io_in_A_2(S8DP1_7_io_in_A_2),
    .io_in_A_3(S8DP1_7_io_in_A_3),
    .io_in_A_4(S8DP1_7_io_in_A_4),
    .io_in_A_5(S8DP1_7_io_in_A_5),
    .io_in_A_6(S8DP1_7_io_in_A_6),
    .io_in_A_7(S8DP1_7_io_in_A_7),
    .io_in_B_0(S8DP1_7_io_in_B_0),
    .io_in_B_1(S8DP1_7_io_in_B_1),
    .io_in_B_2(S8DP1_7_io_in_B_2),
    .io_in_B_3(S8DP1_7_io_in_B_3),
    .io_in_B_4(S8DP1_7_io_in_B_4),
    .io_in_B_5(S8DP1_7_io_in_B_5),
    .io_in_B_6(S8DP1_7_io_in_B_6),
    .io_in_B_7(S8DP1_7_io_in_B_7),
    .io_in_tag_0(S8DP1_7_io_in_tag_0),
    .io_in_tag_1(S8DP1_7_io_in_tag_1),
    .io_in_tag_2(S8DP1_7_io_in_tag_2),
    .io_in_tag_3(S8DP1_7_io_in_tag_3),
    .io_in_tag_4(S8DP1_7_io_in_tag_4),
    .io_in_tag_5(S8DP1_7_io_in_tag_5),
    .io_in_tag_6(S8DP1_7_io_in_tag_6),
    .io_in_tag_7(S8DP1_7_io_in_tag_7),
    .io_result(S8DP1_7_io_result),
    .io_in_calculate(S8DP1_7_io_in_calculate),
    .io_out_calculate(S8DP1_7_io_out_calculate)
  );
  assign S8DP1_1_1_0_out_calculate = S8DP1_io_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1814.4]
  assign S8DP1_1_1_1_out_calculate = S8DP1_1_io_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1841.4]
  assign _T_3683 = S8DP1_1_1_0_out_calculate & S8DP1_1_1_1_out_calculate; // @[TPU.scala 78:42:@2245.4]
  assign S8DP1_1_1_2_out_calculate = S8DP1_2_io_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1868.4]
  assign _T_3684 = _T_3683 & S8DP1_1_1_2_out_calculate; // @[TPU.scala 78:70:@2246.4]
  assign S8DP1_1_1_3_out_calculate = S8DP1_3_io_out_calculate; // @[TPU.scala 62:20:@1813.4 TPU.scala 62:20:@1895.4]
  assign _T_3685 = _T_3684 & S8DP1_1_1_3_out_calculate; // @[TPU.scala 78:98:@2247.4]
  assign S8DP1_2_1_0_out_calculate = S8DP1_4_io_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1935.4]
  assign _T_3686 = _T_3685 & S8DP1_2_1_0_out_calculate; // @[TPU.scala 79:5:@2248.4]
  assign S8DP1_2_1_1_out_calculate = S8DP1_5_io_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1962.4]
  assign _T_3687 = _T_3686 & S8DP1_2_1_1_out_calculate; // @[TPU.scala 79:33:@2249.4]
  assign S8DP1_2_1_2_out_calculate = S8DP1_6_io_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@1989.4]
  assign _T_3688 = _T_3687 & S8DP1_2_1_2_out_calculate; // @[TPU.scala 79:61:@2250.4]
  assign S8DP1_2_1_3_out_calculate = S8DP1_7_io_out_calculate; // @[TPU.scala 63:20:@1934.4 TPU.scala 63:20:@2016.4]
  assign _T_3689 = _T_3688 & S8DP1_2_1_3_out_calculate; // @[TPU.scala 79:89:@2251.4]
  assign _T_3691 = 2'h2 == stateReg; // @[Conditional.scala 37:30:@2263.4]
  assign _T_3695 = _T_3693 == 1'h0; // @[TPU.scala 93:25:@2267.6]
  assign _T_3696 = io_in_cal & _T_3695; // @[TPU.scala 93:23:@2268.6]
  assign _GEN_0 = _T_3696 ? 2'h0 : stateReg; // @[TPU.scala 93:46:@2269.6]
  assign _T_3697 = 2'h0 == stateReg; // @[Conditional.scala 37:30:@2274.6]
  assign _T_3698 = 2'h1 == stateReg; // @[Conditional.scala 37:30:@2279.8]
  assign _GEN_1 = cal_state ? 2'h2 : stateReg; // @[TPU.scala 106:23:@2282.10]
  assign _GEN_2 = cal_state ? 1'h0 : 1'h1; // @[TPU.scala 106:23:@2282.10]
  assign _GEN_3 = _T_3698 ? _GEN_2 : cal_control; // @[Conditional.scala 39:67:@2280.8]
  assign _GEN_4 = _T_3698 ? _GEN_1 : stateReg; // @[Conditional.scala 39:67:@2280.8]
  assign _GEN_5 = _T_3697 ? 2'h1 : _GEN_4; // @[Conditional.scala 39:67:@2275.6]
  assign _GEN_6 = _T_3697 ? cal_control : _GEN_3; // @[Conditional.scala 39:67:@2275.6]
  assign _GEN_7 = _T_3691 ? _GEN_0 : _GEN_5; // @[Conditional.scala 40:58:@2264.4]
  assign _GEN_8 = _T_3691 ? cal_control : _GEN_6; // @[Conditional.scala 40:58:@2264.4]
  assign io_out_A_0_0 = io_in_A_0_0; // @[TPU.scala 54:12:@1721.4]
  assign io_out_A_0_1 = io_in_A_0_1; // @[TPU.scala 54:12:@1722.4]
  assign io_out_A_0_2 = io_in_A_0_2; // @[TPU.scala 54:12:@1723.4]
  assign io_out_A_0_3 = io_in_A_0_3; // @[TPU.scala 54:12:@1724.4]
  assign io_out_A_0_4 = io_in_A_0_4; // @[TPU.scala 54:12:@1725.4]
  assign io_out_A_0_5 = io_in_A_0_5; // @[TPU.scala 54:12:@1726.4]
  assign io_out_A_0_6 = io_in_A_0_6; // @[TPU.scala 54:12:@1727.4]
  assign io_out_A_0_7 = io_in_A_0_7; // @[TPU.scala 54:12:@1728.4]
  assign io_out_A_1_0 = io_in_A_1_0; // @[TPU.scala 54:12:@1729.4]
  assign io_out_A_1_1 = io_in_A_1_1; // @[TPU.scala 54:12:@1730.4]
  assign io_out_A_1_2 = io_in_A_1_2; // @[TPU.scala 54:12:@1731.4]
  assign io_out_A_1_3 = io_in_A_1_3; // @[TPU.scala 54:12:@1732.4]
  assign io_out_A_1_4 = io_in_A_1_4; // @[TPU.scala 54:12:@1733.4]
  assign io_out_A_1_5 = io_in_A_1_5; // @[TPU.scala 54:12:@1734.4]
  assign io_out_A_1_6 = io_in_A_1_6; // @[TPU.scala 54:12:@1735.4]
  assign io_out_A_1_7 = io_in_A_1_7; // @[TPU.scala 54:12:@1736.4]
  assign io_out_B_0_0 = io_in_B_0_0; // @[TPU.scala 57:12:@1737.4]
  assign io_out_B_0_1 = io_in_B_0_1; // @[TPU.scala 57:12:@1738.4]
  assign io_out_B_0_2 = io_in_B_0_2; // @[TPU.scala 57:12:@1739.4]
  assign io_out_B_0_3 = io_in_B_0_3; // @[TPU.scala 57:12:@1740.4]
  assign io_out_B_0_4 = io_in_B_0_4; // @[TPU.scala 57:12:@1741.4]
  assign io_out_B_0_5 = io_in_B_0_5; // @[TPU.scala 57:12:@1742.4]
  assign io_out_B_0_6 = io_in_B_0_6; // @[TPU.scala 57:12:@1743.4]
  assign io_out_B_0_7 = io_in_B_0_7; // @[TPU.scala 57:12:@1744.4]
  assign io_out_B_1_0 = io_in_B_1_0; // @[TPU.scala 57:12:@1745.4]
  assign io_out_B_1_1 = io_in_B_1_1; // @[TPU.scala 57:12:@1746.4]
  assign io_out_B_1_2 = io_in_B_1_2; // @[TPU.scala 57:12:@1747.4]
  assign io_out_B_1_3 = io_in_B_1_3; // @[TPU.scala 57:12:@1748.4]
  assign io_out_B_1_4 = io_in_B_1_4; // @[TPU.scala 57:12:@1749.4]
  assign io_out_B_1_5 = io_in_B_1_5; // @[TPU.scala 57:12:@1750.4]
  assign io_out_B_1_6 = io_in_B_1_6; // @[TPU.scala 57:12:@1751.4]
  assign io_out_B_1_7 = io_in_B_1_7; // @[TPU.scala 57:12:@1752.4]
  assign io_out_B_2_0 = io_in_B_2_0; // @[TPU.scala 57:12:@1753.4]
  assign io_out_B_2_1 = io_in_B_2_1; // @[TPU.scala 57:12:@1754.4]
  assign io_out_B_2_2 = io_in_B_2_2; // @[TPU.scala 57:12:@1755.4]
  assign io_out_B_2_3 = io_in_B_2_3; // @[TPU.scala 57:12:@1756.4]
  assign io_out_B_2_4 = io_in_B_2_4; // @[TPU.scala 57:12:@1757.4]
  assign io_out_B_2_5 = io_in_B_2_5; // @[TPU.scala 57:12:@1758.4]
  assign io_out_B_2_6 = io_in_B_2_6; // @[TPU.scala 57:12:@1759.4]
  assign io_out_B_2_7 = io_in_B_2_7; // @[TPU.scala 57:12:@1760.4]
  assign io_out_B_3_0 = io_in_B_3_0; // @[TPU.scala 57:12:@1761.4]
  assign io_out_B_3_1 = io_in_B_3_1; // @[TPU.scala 57:12:@1762.4]
  assign io_out_B_3_2 = io_in_B_3_2; // @[TPU.scala 57:12:@1763.4]
  assign io_out_B_3_3 = io_in_B_3_3; // @[TPU.scala 57:12:@1764.4]
  assign io_out_B_3_4 = io_in_B_3_4; // @[TPU.scala 57:12:@1765.4]
  assign io_out_B_3_5 = io_in_B_3_5; // @[TPU.scala 57:12:@1766.4]
  assign io_out_B_3_6 = io_in_B_3_6; // @[TPU.scala 57:12:@1767.4]
  assign io_out_B_3_7 = io_in_B_3_7; // @[TPU.scala 57:12:@1768.4]
  assign io_out_tag_0_0 = io_in_tag_0_0; // @[TPU.scala 60:14:@1769.4]
  assign io_out_tag_0_1 = io_in_tag_0_1; // @[TPU.scala 60:14:@1770.4]
  assign io_out_tag_0_2 = io_in_tag_0_2; // @[TPU.scala 60:14:@1771.4]
  assign io_out_tag_0_3 = io_in_tag_0_3; // @[TPU.scala 60:14:@1772.4]
  assign io_out_tag_0_4 = io_in_tag_0_4; // @[TPU.scala 60:14:@1773.4]
  assign io_out_tag_0_5 = io_in_tag_0_5; // @[TPU.scala 60:14:@1774.4]
  assign io_out_tag_0_6 = io_in_tag_0_6; // @[TPU.scala 60:14:@1775.4]
  assign io_out_tag_0_7 = io_in_tag_0_7; // @[TPU.scala 60:14:@1776.4]
  assign io_out_tag_1_0 = io_in_tag_1_0; // @[TPU.scala 60:14:@1777.4]
  assign io_out_tag_1_1 = io_in_tag_1_1; // @[TPU.scala 60:14:@1778.4]
  assign io_out_tag_1_2 = io_in_tag_1_2; // @[TPU.scala 60:14:@1779.4]
  assign io_out_tag_1_3 = io_in_tag_1_3; // @[TPU.scala 60:14:@1780.4]
  assign io_out_tag_1_4 = io_in_tag_1_4; // @[TPU.scala 60:14:@1781.4]
  assign io_out_tag_1_5 = io_in_tag_1_5; // @[TPU.scala 60:14:@1782.4]
  assign io_out_tag_1_6 = io_in_tag_1_6; // @[TPU.scala 60:14:@1783.4]
  assign io_out_tag_1_7 = io_in_tag_1_7; // @[TPU.scala 60:14:@1784.4]
  assign io_out_tag_2_0 = io_in_tag_2_0; // @[TPU.scala 60:14:@1785.4]
  assign io_out_tag_2_1 = io_in_tag_2_1; // @[TPU.scala 60:14:@1786.4]
  assign io_out_tag_2_2 = io_in_tag_2_2; // @[TPU.scala 60:14:@1787.4]
  assign io_out_tag_2_3 = io_in_tag_2_3; // @[TPU.scala 60:14:@1788.4]
  assign io_out_tag_2_4 = io_in_tag_2_4; // @[TPU.scala 60:14:@1789.4]
  assign io_out_tag_2_5 = io_in_tag_2_5; // @[TPU.scala 60:14:@1790.4]
  assign io_out_tag_2_6 = io_in_tag_2_6; // @[TPU.scala 60:14:@1791.4]
  assign io_out_tag_2_7 = io_in_tag_2_7; // @[TPU.scala 60:14:@1792.4]
  assign io_out_tag_3_0 = io_in_tag_3_0; // @[TPU.scala 60:14:@1793.4]
  assign io_out_tag_3_1 = io_in_tag_3_1; // @[TPU.scala 60:14:@1794.4]
  assign io_out_tag_3_2 = io_in_tag_3_2; // @[TPU.scala 60:14:@1795.4]
  assign io_out_tag_3_3 = io_in_tag_3_3; // @[TPU.scala 60:14:@1796.4]
  assign io_out_tag_3_4 = io_in_tag_3_4; // @[TPU.scala 60:14:@1797.4]
  assign io_out_tag_3_5 = io_in_tag_3_5; // @[TPU.scala 60:14:@1798.4]
  assign io_out_tag_3_6 = io_in_tag_3_6; // @[TPU.scala 60:14:@1799.4]
  assign io_out_tag_3_7 = io_in_tag_3_7; // @[TPU.scala 60:14:@1800.4]
  assign io_out_result_0_0 = S8DP1_io_result; // @[TPU.scala 83:25:@2253.4]
  assign io_out_result_0_1 = S8DP1_1_io_result; // @[TPU.scala 83:25:@2255.4]
  assign io_out_result_0_2 = S8DP1_2_io_result; // @[TPU.scala 83:25:@2257.4]
  assign io_out_result_0_3 = S8DP1_3_io_result; // @[TPU.scala 83:25:@2259.4]
  assign io_out_result_1_0 = S8DP1_4_io_result; // @[TPU.scala 84:25:@2254.4]
  assign io_out_result_1_1 = S8DP1_5_io_result; // @[TPU.scala 84:25:@2256.4]
  assign io_out_result_1_2 = S8DP1_6_io_result; // @[TPU.scala 84:25:@2258.4]
  assign io_out_result_1_3 = S8DP1_7_io_result; // @[TPU.scala 84:25:@2260.4]
  assign io_out_cal = cal_state; // @[TPU.scala 86:14:@2261.4]
  assign S8DP1_clock = clock; // @[:@1802.4]
  assign S8DP1_reset = reset; // @[:@1803.4]
  assign S8DP1_io_in_A_0 = io_in_A_0_0; // @[TPU.scala 62:20:@1833.4]
  assign S8DP1_io_in_A_1 = io_in_A_0_1; // @[TPU.scala 62:20:@1834.4]
  assign S8DP1_io_in_A_2 = io_in_A_0_2; // @[TPU.scala 62:20:@1835.4]
  assign S8DP1_io_in_A_3 = io_in_A_0_3; // @[TPU.scala 62:20:@1836.4]
  assign S8DP1_io_in_A_4 = io_in_A_0_4; // @[TPU.scala 62:20:@1837.4]
  assign S8DP1_io_in_A_5 = io_in_A_0_5; // @[TPU.scala 62:20:@1838.4]
  assign S8DP1_io_in_A_6 = io_in_A_0_6; // @[TPU.scala 62:20:@1839.4]
  assign S8DP1_io_in_A_7 = io_in_A_0_7; // @[TPU.scala 62:20:@1840.4]
  assign S8DP1_io_in_B_0 = io_in_B_0_0; // @[TPU.scala 62:20:@1825.4]
  assign S8DP1_io_in_B_1 = io_in_B_0_1; // @[TPU.scala 62:20:@1826.4]
  assign S8DP1_io_in_B_2 = io_in_B_0_2; // @[TPU.scala 62:20:@1827.4]
  assign S8DP1_io_in_B_3 = io_in_B_0_3; // @[TPU.scala 62:20:@1828.4]
  assign S8DP1_io_in_B_4 = io_in_B_0_4; // @[TPU.scala 62:20:@1829.4]
  assign S8DP1_io_in_B_5 = io_in_B_0_5; // @[TPU.scala 62:20:@1830.4]
  assign S8DP1_io_in_B_6 = io_in_B_0_6; // @[TPU.scala 62:20:@1831.4]
  assign S8DP1_io_in_B_7 = io_in_B_0_7; // @[TPU.scala 62:20:@1832.4]
  assign S8DP1_io_in_tag_0 = io_in_tag_0_0; // @[TPU.scala 62:20:@1817.4]
  assign S8DP1_io_in_tag_1 = io_in_tag_0_1; // @[TPU.scala 62:20:@1818.4]
  assign S8DP1_io_in_tag_2 = io_in_tag_0_2; // @[TPU.scala 62:20:@1819.4]
  assign S8DP1_io_in_tag_3 = io_in_tag_0_3; // @[TPU.scala 62:20:@1820.4]
  assign S8DP1_io_in_tag_4 = io_in_tag_0_4; // @[TPU.scala 62:20:@1821.4]
  assign S8DP1_io_in_tag_5 = io_in_tag_0_5; // @[TPU.scala 62:20:@1822.4]
  assign S8DP1_io_in_tag_6 = io_in_tag_0_6; // @[TPU.scala 62:20:@1823.4]
  assign S8DP1_io_in_tag_7 = io_in_tag_0_7; // @[TPU.scala 62:20:@1824.4]
  assign S8DP1_io_in_calculate = cal_control; // @[TPU.scala 62:20:@1815.4]
  assign S8DP1_1_clock = clock; // @[:@1805.4]
  assign S8DP1_1_reset = reset; // @[:@1806.4]
  assign S8DP1_1_io_in_A_0 = io_in_A_0_0; // @[TPU.scala 62:20:@1860.4]
  assign S8DP1_1_io_in_A_1 = io_in_A_0_1; // @[TPU.scala 62:20:@1861.4]
  assign S8DP1_1_io_in_A_2 = io_in_A_0_2; // @[TPU.scala 62:20:@1862.4]
  assign S8DP1_1_io_in_A_3 = io_in_A_0_3; // @[TPU.scala 62:20:@1863.4]
  assign S8DP1_1_io_in_A_4 = io_in_A_0_4; // @[TPU.scala 62:20:@1864.4]
  assign S8DP1_1_io_in_A_5 = io_in_A_0_5; // @[TPU.scala 62:20:@1865.4]
  assign S8DP1_1_io_in_A_6 = io_in_A_0_6; // @[TPU.scala 62:20:@1866.4]
  assign S8DP1_1_io_in_A_7 = io_in_A_0_7; // @[TPU.scala 62:20:@1867.4]
  assign S8DP1_1_io_in_B_0 = io_in_B_1_0; // @[TPU.scala 62:20:@1852.4]
  assign S8DP1_1_io_in_B_1 = io_in_B_1_1; // @[TPU.scala 62:20:@1853.4]
  assign S8DP1_1_io_in_B_2 = io_in_B_1_2; // @[TPU.scala 62:20:@1854.4]
  assign S8DP1_1_io_in_B_3 = io_in_B_1_3; // @[TPU.scala 62:20:@1855.4]
  assign S8DP1_1_io_in_B_4 = io_in_B_1_4; // @[TPU.scala 62:20:@1856.4]
  assign S8DP1_1_io_in_B_5 = io_in_B_1_5; // @[TPU.scala 62:20:@1857.4]
  assign S8DP1_1_io_in_B_6 = io_in_B_1_6; // @[TPU.scala 62:20:@1858.4]
  assign S8DP1_1_io_in_B_7 = io_in_B_1_7; // @[TPU.scala 62:20:@1859.4]
  assign S8DP1_1_io_in_tag_0 = io_in_tag_1_0; // @[TPU.scala 62:20:@1844.4]
  assign S8DP1_1_io_in_tag_1 = io_in_tag_1_1; // @[TPU.scala 62:20:@1845.4]
  assign S8DP1_1_io_in_tag_2 = io_in_tag_1_2; // @[TPU.scala 62:20:@1846.4]
  assign S8DP1_1_io_in_tag_3 = io_in_tag_1_3; // @[TPU.scala 62:20:@1847.4]
  assign S8DP1_1_io_in_tag_4 = io_in_tag_1_4; // @[TPU.scala 62:20:@1848.4]
  assign S8DP1_1_io_in_tag_5 = io_in_tag_1_5; // @[TPU.scala 62:20:@1849.4]
  assign S8DP1_1_io_in_tag_6 = io_in_tag_1_6; // @[TPU.scala 62:20:@1850.4]
  assign S8DP1_1_io_in_tag_7 = io_in_tag_1_7; // @[TPU.scala 62:20:@1851.4]
  assign S8DP1_1_io_in_calculate = cal_control; // @[TPU.scala 62:20:@1842.4]
  assign S8DP1_2_clock = clock; // @[:@1808.4]
  assign S8DP1_2_reset = reset; // @[:@1809.4]
  assign S8DP1_2_io_in_A_0 = io_in_A_0_0; // @[TPU.scala 62:20:@1887.4]
  assign S8DP1_2_io_in_A_1 = io_in_A_0_1; // @[TPU.scala 62:20:@1888.4]
  assign S8DP1_2_io_in_A_2 = io_in_A_0_2; // @[TPU.scala 62:20:@1889.4]
  assign S8DP1_2_io_in_A_3 = io_in_A_0_3; // @[TPU.scala 62:20:@1890.4]
  assign S8DP1_2_io_in_A_4 = io_in_A_0_4; // @[TPU.scala 62:20:@1891.4]
  assign S8DP1_2_io_in_A_5 = io_in_A_0_5; // @[TPU.scala 62:20:@1892.4]
  assign S8DP1_2_io_in_A_6 = io_in_A_0_6; // @[TPU.scala 62:20:@1893.4]
  assign S8DP1_2_io_in_A_7 = io_in_A_0_7; // @[TPU.scala 62:20:@1894.4]
  assign S8DP1_2_io_in_B_0 = io_in_B_2_0; // @[TPU.scala 62:20:@1879.4]
  assign S8DP1_2_io_in_B_1 = io_in_B_2_1; // @[TPU.scala 62:20:@1880.4]
  assign S8DP1_2_io_in_B_2 = io_in_B_2_2; // @[TPU.scala 62:20:@1881.4]
  assign S8DP1_2_io_in_B_3 = io_in_B_2_3; // @[TPU.scala 62:20:@1882.4]
  assign S8DP1_2_io_in_B_4 = io_in_B_2_4; // @[TPU.scala 62:20:@1883.4]
  assign S8DP1_2_io_in_B_5 = io_in_B_2_5; // @[TPU.scala 62:20:@1884.4]
  assign S8DP1_2_io_in_B_6 = io_in_B_2_6; // @[TPU.scala 62:20:@1885.4]
  assign S8DP1_2_io_in_B_7 = io_in_B_2_7; // @[TPU.scala 62:20:@1886.4]
  assign S8DP1_2_io_in_tag_0 = io_in_tag_2_0; // @[TPU.scala 62:20:@1871.4]
  assign S8DP1_2_io_in_tag_1 = io_in_tag_2_1; // @[TPU.scala 62:20:@1872.4]
  assign S8DP1_2_io_in_tag_2 = io_in_tag_2_2; // @[TPU.scala 62:20:@1873.4]
  assign S8DP1_2_io_in_tag_3 = io_in_tag_2_3; // @[TPU.scala 62:20:@1874.4]
  assign S8DP1_2_io_in_tag_4 = io_in_tag_2_4; // @[TPU.scala 62:20:@1875.4]
  assign S8DP1_2_io_in_tag_5 = io_in_tag_2_5; // @[TPU.scala 62:20:@1876.4]
  assign S8DP1_2_io_in_tag_6 = io_in_tag_2_6; // @[TPU.scala 62:20:@1877.4]
  assign S8DP1_2_io_in_tag_7 = io_in_tag_2_7; // @[TPU.scala 62:20:@1878.4]
  assign S8DP1_2_io_in_calculate = cal_control; // @[TPU.scala 62:20:@1869.4]
  assign S8DP1_3_clock = clock; // @[:@1811.4]
  assign S8DP1_3_reset = reset; // @[:@1812.4]
  assign S8DP1_3_io_in_A_0 = io_in_A_0_0; // @[TPU.scala 62:20:@1914.4]
  assign S8DP1_3_io_in_A_1 = io_in_A_0_1; // @[TPU.scala 62:20:@1915.4]
  assign S8DP1_3_io_in_A_2 = io_in_A_0_2; // @[TPU.scala 62:20:@1916.4]
  assign S8DP1_3_io_in_A_3 = io_in_A_0_3; // @[TPU.scala 62:20:@1917.4]
  assign S8DP1_3_io_in_A_4 = io_in_A_0_4; // @[TPU.scala 62:20:@1918.4]
  assign S8DP1_3_io_in_A_5 = io_in_A_0_5; // @[TPU.scala 62:20:@1919.4]
  assign S8DP1_3_io_in_A_6 = io_in_A_0_6; // @[TPU.scala 62:20:@1920.4]
  assign S8DP1_3_io_in_A_7 = io_in_A_0_7; // @[TPU.scala 62:20:@1921.4]
  assign S8DP1_3_io_in_B_0 = io_in_B_3_0; // @[TPU.scala 62:20:@1906.4]
  assign S8DP1_3_io_in_B_1 = io_in_B_3_1; // @[TPU.scala 62:20:@1907.4]
  assign S8DP1_3_io_in_B_2 = io_in_B_3_2; // @[TPU.scala 62:20:@1908.4]
  assign S8DP1_3_io_in_B_3 = io_in_B_3_3; // @[TPU.scala 62:20:@1909.4]
  assign S8DP1_3_io_in_B_4 = io_in_B_3_4; // @[TPU.scala 62:20:@1910.4]
  assign S8DP1_3_io_in_B_5 = io_in_B_3_5; // @[TPU.scala 62:20:@1911.4]
  assign S8DP1_3_io_in_B_6 = io_in_B_3_6; // @[TPU.scala 62:20:@1912.4]
  assign S8DP1_3_io_in_B_7 = io_in_B_3_7; // @[TPU.scala 62:20:@1913.4]
  assign S8DP1_3_io_in_tag_0 = io_in_tag_3_0; // @[TPU.scala 62:20:@1898.4]
  assign S8DP1_3_io_in_tag_1 = io_in_tag_3_1; // @[TPU.scala 62:20:@1899.4]
  assign S8DP1_3_io_in_tag_2 = io_in_tag_3_2; // @[TPU.scala 62:20:@1900.4]
  assign S8DP1_3_io_in_tag_3 = io_in_tag_3_3; // @[TPU.scala 62:20:@1901.4]
  assign S8DP1_3_io_in_tag_4 = io_in_tag_3_4; // @[TPU.scala 62:20:@1902.4]
  assign S8DP1_3_io_in_tag_5 = io_in_tag_3_5; // @[TPU.scala 62:20:@1903.4]
  assign S8DP1_3_io_in_tag_6 = io_in_tag_3_6; // @[TPU.scala 62:20:@1904.4]
  assign S8DP1_3_io_in_tag_7 = io_in_tag_3_7; // @[TPU.scala 62:20:@1905.4]
  assign S8DP1_3_io_in_calculate = cal_control; // @[TPU.scala 62:20:@1896.4]
  assign S8DP1_4_clock = clock; // @[:@1923.4]
  assign S8DP1_4_reset = reset; // @[:@1924.4]
  assign S8DP1_4_io_in_A_0 = io_in_A_1_0; // @[TPU.scala 63:20:@1954.4]
  assign S8DP1_4_io_in_A_1 = io_in_A_1_1; // @[TPU.scala 63:20:@1955.4]
  assign S8DP1_4_io_in_A_2 = io_in_A_1_2; // @[TPU.scala 63:20:@1956.4]
  assign S8DP1_4_io_in_A_3 = io_in_A_1_3; // @[TPU.scala 63:20:@1957.4]
  assign S8DP1_4_io_in_A_4 = io_in_A_1_4; // @[TPU.scala 63:20:@1958.4]
  assign S8DP1_4_io_in_A_5 = io_in_A_1_5; // @[TPU.scala 63:20:@1959.4]
  assign S8DP1_4_io_in_A_6 = io_in_A_1_6; // @[TPU.scala 63:20:@1960.4]
  assign S8DP1_4_io_in_A_7 = io_in_A_1_7; // @[TPU.scala 63:20:@1961.4]
  assign S8DP1_4_io_in_B_0 = io_in_B_0_0; // @[TPU.scala 63:20:@1946.4]
  assign S8DP1_4_io_in_B_1 = io_in_B_0_1; // @[TPU.scala 63:20:@1947.4]
  assign S8DP1_4_io_in_B_2 = io_in_B_0_2; // @[TPU.scala 63:20:@1948.4]
  assign S8DP1_4_io_in_B_3 = io_in_B_0_3; // @[TPU.scala 63:20:@1949.4]
  assign S8DP1_4_io_in_B_4 = io_in_B_0_4; // @[TPU.scala 63:20:@1950.4]
  assign S8DP1_4_io_in_B_5 = io_in_B_0_5; // @[TPU.scala 63:20:@1951.4]
  assign S8DP1_4_io_in_B_6 = io_in_B_0_6; // @[TPU.scala 63:20:@1952.4]
  assign S8DP1_4_io_in_B_7 = io_in_B_0_7; // @[TPU.scala 63:20:@1953.4]
  assign S8DP1_4_io_in_tag_0 = io_in_tag_0_0; // @[TPU.scala 63:20:@1938.4]
  assign S8DP1_4_io_in_tag_1 = io_in_tag_0_1; // @[TPU.scala 63:20:@1939.4]
  assign S8DP1_4_io_in_tag_2 = io_in_tag_0_2; // @[TPU.scala 63:20:@1940.4]
  assign S8DP1_4_io_in_tag_3 = io_in_tag_0_3; // @[TPU.scala 63:20:@1941.4]
  assign S8DP1_4_io_in_tag_4 = io_in_tag_0_4; // @[TPU.scala 63:20:@1942.4]
  assign S8DP1_4_io_in_tag_5 = io_in_tag_0_5; // @[TPU.scala 63:20:@1943.4]
  assign S8DP1_4_io_in_tag_6 = io_in_tag_0_6; // @[TPU.scala 63:20:@1944.4]
  assign S8DP1_4_io_in_tag_7 = io_in_tag_0_7; // @[TPU.scala 63:20:@1945.4]
  assign S8DP1_4_io_in_calculate = cal_control; // @[TPU.scala 63:20:@1936.4]
  assign S8DP1_5_clock = clock; // @[:@1926.4]
  assign S8DP1_5_reset = reset; // @[:@1927.4]
  assign S8DP1_5_io_in_A_0 = io_in_A_1_0; // @[TPU.scala 63:20:@1981.4]
  assign S8DP1_5_io_in_A_1 = io_in_A_1_1; // @[TPU.scala 63:20:@1982.4]
  assign S8DP1_5_io_in_A_2 = io_in_A_1_2; // @[TPU.scala 63:20:@1983.4]
  assign S8DP1_5_io_in_A_3 = io_in_A_1_3; // @[TPU.scala 63:20:@1984.4]
  assign S8DP1_5_io_in_A_4 = io_in_A_1_4; // @[TPU.scala 63:20:@1985.4]
  assign S8DP1_5_io_in_A_5 = io_in_A_1_5; // @[TPU.scala 63:20:@1986.4]
  assign S8DP1_5_io_in_A_6 = io_in_A_1_6; // @[TPU.scala 63:20:@1987.4]
  assign S8DP1_5_io_in_A_7 = io_in_A_1_7; // @[TPU.scala 63:20:@1988.4]
  assign S8DP1_5_io_in_B_0 = io_in_B_1_0; // @[TPU.scala 63:20:@1973.4]
  assign S8DP1_5_io_in_B_1 = io_in_B_1_1; // @[TPU.scala 63:20:@1974.4]
  assign S8DP1_5_io_in_B_2 = io_in_B_1_2; // @[TPU.scala 63:20:@1975.4]
  assign S8DP1_5_io_in_B_3 = io_in_B_1_3; // @[TPU.scala 63:20:@1976.4]
  assign S8DP1_5_io_in_B_4 = io_in_B_1_4; // @[TPU.scala 63:20:@1977.4]
  assign S8DP1_5_io_in_B_5 = io_in_B_1_5; // @[TPU.scala 63:20:@1978.4]
  assign S8DP1_5_io_in_B_6 = io_in_B_1_6; // @[TPU.scala 63:20:@1979.4]
  assign S8DP1_5_io_in_B_7 = io_in_B_1_7; // @[TPU.scala 63:20:@1980.4]
  assign S8DP1_5_io_in_tag_0 = io_in_tag_1_0; // @[TPU.scala 63:20:@1965.4]
  assign S8DP1_5_io_in_tag_1 = io_in_tag_1_1; // @[TPU.scala 63:20:@1966.4]
  assign S8DP1_5_io_in_tag_2 = io_in_tag_1_2; // @[TPU.scala 63:20:@1967.4]
  assign S8DP1_5_io_in_tag_3 = io_in_tag_1_3; // @[TPU.scala 63:20:@1968.4]
  assign S8DP1_5_io_in_tag_4 = io_in_tag_1_4; // @[TPU.scala 63:20:@1969.4]
  assign S8DP1_5_io_in_tag_5 = io_in_tag_1_5; // @[TPU.scala 63:20:@1970.4]
  assign S8DP1_5_io_in_tag_6 = io_in_tag_1_6; // @[TPU.scala 63:20:@1971.4]
  assign S8DP1_5_io_in_tag_7 = io_in_tag_1_7; // @[TPU.scala 63:20:@1972.4]
  assign S8DP1_5_io_in_calculate = cal_control; // @[TPU.scala 63:20:@1963.4]
  assign S8DP1_6_clock = clock; // @[:@1929.4]
  assign S8DP1_6_reset = reset; // @[:@1930.4]
  assign S8DP1_6_io_in_A_0 = io_in_A_1_0; // @[TPU.scala 63:20:@2008.4]
  assign S8DP1_6_io_in_A_1 = io_in_A_1_1; // @[TPU.scala 63:20:@2009.4]
  assign S8DP1_6_io_in_A_2 = io_in_A_1_2; // @[TPU.scala 63:20:@2010.4]
  assign S8DP1_6_io_in_A_3 = io_in_A_1_3; // @[TPU.scala 63:20:@2011.4]
  assign S8DP1_6_io_in_A_4 = io_in_A_1_4; // @[TPU.scala 63:20:@2012.4]
  assign S8DP1_6_io_in_A_5 = io_in_A_1_5; // @[TPU.scala 63:20:@2013.4]
  assign S8DP1_6_io_in_A_6 = io_in_A_1_6; // @[TPU.scala 63:20:@2014.4]
  assign S8DP1_6_io_in_A_7 = io_in_A_1_7; // @[TPU.scala 63:20:@2015.4]
  assign S8DP1_6_io_in_B_0 = io_in_B_2_0; // @[TPU.scala 63:20:@2000.4]
  assign S8DP1_6_io_in_B_1 = io_in_B_2_1; // @[TPU.scala 63:20:@2001.4]
  assign S8DP1_6_io_in_B_2 = io_in_B_2_2; // @[TPU.scala 63:20:@2002.4]
  assign S8DP1_6_io_in_B_3 = io_in_B_2_3; // @[TPU.scala 63:20:@2003.4]
  assign S8DP1_6_io_in_B_4 = io_in_B_2_4; // @[TPU.scala 63:20:@2004.4]
  assign S8DP1_6_io_in_B_5 = io_in_B_2_5; // @[TPU.scala 63:20:@2005.4]
  assign S8DP1_6_io_in_B_6 = io_in_B_2_6; // @[TPU.scala 63:20:@2006.4]
  assign S8DP1_6_io_in_B_7 = io_in_B_2_7; // @[TPU.scala 63:20:@2007.4]
  assign S8DP1_6_io_in_tag_0 = io_in_tag_2_0; // @[TPU.scala 63:20:@1992.4]
  assign S8DP1_6_io_in_tag_1 = io_in_tag_2_1; // @[TPU.scala 63:20:@1993.4]
  assign S8DP1_6_io_in_tag_2 = io_in_tag_2_2; // @[TPU.scala 63:20:@1994.4]
  assign S8DP1_6_io_in_tag_3 = io_in_tag_2_3; // @[TPU.scala 63:20:@1995.4]
  assign S8DP1_6_io_in_tag_4 = io_in_tag_2_4; // @[TPU.scala 63:20:@1996.4]
  assign S8DP1_6_io_in_tag_5 = io_in_tag_2_5; // @[TPU.scala 63:20:@1997.4]
  assign S8DP1_6_io_in_tag_6 = io_in_tag_2_6; // @[TPU.scala 63:20:@1998.4]
  assign S8DP1_6_io_in_tag_7 = io_in_tag_2_7; // @[TPU.scala 63:20:@1999.4]
  assign S8DP1_6_io_in_calculate = cal_control; // @[TPU.scala 63:20:@1990.4]
  assign S8DP1_7_clock = clock; // @[:@1932.4]
  assign S8DP1_7_reset = reset; // @[:@1933.4]
  assign S8DP1_7_io_in_A_0 = io_in_A_1_0; // @[TPU.scala 63:20:@2035.4]
  assign S8DP1_7_io_in_A_1 = io_in_A_1_1; // @[TPU.scala 63:20:@2036.4]
  assign S8DP1_7_io_in_A_2 = io_in_A_1_2; // @[TPU.scala 63:20:@2037.4]
  assign S8DP1_7_io_in_A_3 = io_in_A_1_3; // @[TPU.scala 63:20:@2038.4]
  assign S8DP1_7_io_in_A_4 = io_in_A_1_4; // @[TPU.scala 63:20:@2039.4]
  assign S8DP1_7_io_in_A_5 = io_in_A_1_5; // @[TPU.scala 63:20:@2040.4]
  assign S8DP1_7_io_in_A_6 = io_in_A_1_6; // @[TPU.scala 63:20:@2041.4]
  assign S8DP1_7_io_in_A_7 = io_in_A_1_7; // @[TPU.scala 63:20:@2042.4]
  assign S8DP1_7_io_in_B_0 = io_in_B_3_0; // @[TPU.scala 63:20:@2027.4]
  assign S8DP1_7_io_in_B_1 = io_in_B_3_1; // @[TPU.scala 63:20:@2028.4]
  assign S8DP1_7_io_in_B_2 = io_in_B_3_2; // @[TPU.scala 63:20:@2029.4]
  assign S8DP1_7_io_in_B_3 = io_in_B_3_3; // @[TPU.scala 63:20:@2030.4]
  assign S8DP1_7_io_in_B_4 = io_in_B_3_4; // @[TPU.scala 63:20:@2031.4]
  assign S8DP1_7_io_in_B_5 = io_in_B_3_5; // @[TPU.scala 63:20:@2032.4]
  assign S8DP1_7_io_in_B_6 = io_in_B_3_6; // @[TPU.scala 63:20:@2033.4]
  assign S8DP1_7_io_in_B_7 = io_in_B_3_7; // @[TPU.scala 63:20:@2034.4]
  assign S8DP1_7_io_in_tag_0 = io_in_tag_3_0; // @[TPU.scala 63:20:@2019.4]
  assign S8DP1_7_io_in_tag_1 = io_in_tag_3_1; // @[TPU.scala 63:20:@2020.4]
  assign S8DP1_7_io_in_tag_2 = io_in_tag_3_2; // @[TPU.scala 63:20:@2021.4]
  assign S8DP1_7_io_in_tag_3 = io_in_tag_3_3; // @[TPU.scala 63:20:@2022.4]
  assign S8DP1_7_io_in_tag_4 = io_in_tag_3_4; // @[TPU.scala 63:20:@2023.4]
  assign S8DP1_7_io_in_tag_5 = io_in_tag_3_5; // @[TPU.scala 63:20:@2024.4]
  assign S8DP1_7_io_in_tag_6 = io_in_tag_3_6; // @[TPU.scala 63:20:@2025.4]
  assign S8DP1_7_io_in_tag_7 = io_in_tag_3_7; // @[TPU.scala 63:20:@2026.4]
  assign S8DP1_7_io_in_calculate = cal_control; // @[TPU.scala 63:20:@2017.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  cal_state = _RAND_0[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  cal_control = _RAND_1[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  stateReg = _RAND_2[1:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  _T_3693 = _RAND_3[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      cal_state <= 1'h0;
    end else begin
      cal_state <= _T_3689;
    end
    if (reset) begin
      cal_control <= 1'h0;
    end else begin
      if (!(_T_3691)) begin
        if (!(_T_3697)) begin
          if (_T_3698) begin
            if (cal_state) begin
              cal_control <= 1'h0;
            end else begin
              cal_control <= 1'h1;
            end
          end
        end
      end
    end
    if (reset) begin
      stateReg <= 2'h2;
    end else begin
      if (_T_3691) begin
        if (_T_3696) begin
          stateReg <= 2'h0;
        end
      end else begin
        if (_T_3697) begin
          stateReg <= 2'h1;
        end else begin
          if (_T_3698) begin
            if (cal_state) begin
              stateReg <= 2'h2;
            end
          end
        end
      end
    end
    _T_3693 <= io_in_cal;
  end
endmodule
module STA_VDBB( // @[:@7772.2]
  input         clock, // @[:@7773.4]
  input         reset, // @[:@7774.4]
  input  [31:0] io_in_A_0_0, // @[:@7775.4]
  input  [31:0] io_in_A_0_1, // @[:@7775.4]
  input  [31:0] io_in_A_0_2, // @[:@7775.4]
  input  [31:0] io_in_A_0_3, // @[:@7775.4]
  input  [31:0] io_in_A_0_4, // @[:@7775.4]
  input  [31:0] io_in_A_0_5, // @[:@7775.4]
  input  [31:0] io_in_A_0_6, // @[:@7775.4]
  input  [31:0] io_in_A_0_7, // @[:@7775.4]
  input  [31:0] io_in_A_0_8, // @[:@7775.4]
  input  [31:0] io_in_A_0_9, // @[:@7775.4]
  input  [31:0] io_in_A_0_10, // @[:@7775.4]
  input  [31:0] io_in_A_0_11, // @[:@7775.4]
  input  [31:0] io_in_A_0_12, // @[:@7775.4]
  input  [31:0] io_in_A_0_13, // @[:@7775.4]
  input  [31:0] io_in_A_0_14, // @[:@7775.4]
  input  [31:0] io_in_A_0_15, // @[:@7775.4]
  input  [31:0] io_in_A_1_0, // @[:@7775.4]
  input  [31:0] io_in_A_1_1, // @[:@7775.4]
  input  [31:0] io_in_A_1_2, // @[:@7775.4]
  input  [31:0] io_in_A_1_3, // @[:@7775.4]
  input  [31:0] io_in_A_1_4, // @[:@7775.4]
  input  [31:0] io_in_A_1_5, // @[:@7775.4]
  input  [31:0] io_in_A_1_6, // @[:@7775.4]
  input  [31:0] io_in_A_1_7, // @[:@7775.4]
  input  [31:0] io_in_A_1_8, // @[:@7775.4]
  input  [31:0] io_in_A_1_9, // @[:@7775.4]
  input  [31:0] io_in_A_1_10, // @[:@7775.4]
  input  [31:0] io_in_A_1_11, // @[:@7775.4]
  input  [31:0] io_in_A_1_12, // @[:@7775.4]
  input  [31:0] io_in_A_1_13, // @[:@7775.4]
  input  [31:0] io_in_A_1_14, // @[:@7775.4]
  input  [31:0] io_in_A_1_15, // @[:@7775.4]
  input  [31:0] io_in_A_2_0, // @[:@7775.4]
  input  [31:0] io_in_A_2_1, // @[:@7775.4]
  input  [31:0] io_in_A_2_2, // @[:@7775.4]
  input  [31:0] io_in_A_2_3, // @[:@7775.4]
  input  [31:0] io_in_A_2_4, // @[:@7775.4]
  input  [31:0] io_in_A_2_5, // @[:@7775.4]
  input  [31:0] io_in_A_2_6, // @[:@7775.4]
  input  [31:0] io_in_A_2_7, // @[:@7775.4]
  input  [31:0] io_in_A_2_8, // @[:@7775.4]
  input  [31:0] io_in_A_2_9, // @[:@7775.4]
  input  [31:0] io_in_A_2_10, // @[:@7775.4]
  input  [31:0] io_in_A_2_11, // @[:@7775.4]
  input  [31:0] io_in_A_2_12, // @[:@7775.4]
  input  [31:0] io_in_A_2_13, // @[:@7775.4]
  input  [31:0] io_in_A_2_14, // @[:@7775.4]
  input  [31:0] io_in_A_2_15, // @[:@7775.4]
  input  [31:0] io_in_A_3_0, // @[:@7775.4]
  input  [31:0] io_in_A_3_1, // @[:@7775.4]
  input  [31:0] io_in_A_3_2, // @[:@7775.4]
  input  [31:0] io_in_A_3_3, // @[:@7775.4]
  input  [31:0] io_in_A_3_4, // @[:@7775.4]
  input  [31:0] io_in_A_3_5, // @[:@7775.4]
  input  [31:0] io_in_A_3_6, // @[:@7775.4]
  input  [31:0] io_in_A_3_7, // @[:@7775.4]
  input  [31:0] io_in_A_3_8, // @[:@7775.4]
  input  [31:0] io_in_A_3_9, // @[:@7775.4]
  input  [31:0] io_in_A_3_10, // @[:@7775.4]
  input  [31:0] io_in_A_3_11, // @[:@7775.4]
  input  [31:0] io_in_A_3_12, // @[:@7775.4]
  input  [31:0] io_in_A_3_13, // @[:@7775.4]
  input  [31:0] io_in_A_3_14, // @[:@7775.4]
  input  [31:0] io_in_A_3_15, // @[:@7775.4]
  input  [31:0] io_in_B_0_0, // @[:@7775.4]
  input  [31:0] io_in_B_0_1, // @[:@7775.4]
  input  [31:0] io_in_B_0_2, // @[:@7775.4]
  input  [31:0] io_in_B_0_3, // @[:@7775.4]
  input  [31:0] io_in_B_0_4, // @[:@7775.4]
  input  [31:0] io_in_B_0_5, // @[:@7775.4]
  input  [31:0] io_in_B_0_6, // @[:@7775.4]
  input  [31:0] io_in_B_0_7, // @[:@7775.4]
  input  [31:0] io_in_B_0_8, // @[:@7775.4]
  input  [31:0] io_in_B_0_9, // @[:@7775.4]
  input  [31:0] io_in_B_0_10, // @[:@7775.4]
  input  [31:0] io_in_B_0_11, // @[:@7775.4]
  input  [31:0] io_in_B_0_12, // @[:@7775.4]
  input  [31:0] io_in_B_0_13, // @[:@7775.4]
  input  [31:0] io_in_B_0_14, // @[:@7775.4]
  input  [31:0] io_in_B_0_15, // @[:@7775.4]
  input  [31:0] io_in_B_1_0, // @[:@7775.4]
  input  [31:0] io_in_B_1_1, // @[:@7775.4]
  input  [31:0] io_in_B_1_2, // @[:@7775.4]
  input  [31:0] io_in_B_1_3, // @[:@7775.4]
  input  [31:0] io_in_B_1_4, // @[:@7775.4]
  input  [31:0] io_in_B_1_5, // @[:@7775.4]
  input  [31:0] io_in_B_1_6, // @[:@7775.4]
  input  [31:0] io_in_B_1_7, // @[:@7775.4]
  input  [31:0] io_in_B_1_8, // @[:@7775.4]
  input  [31:0] io_in_B_1_9, // @[:@7775.4]
  input  [31:0] io_in_B_1_10, // @[:@7775.4]
  input  [31:0] io_in_B_1_11, // @[:@7775.4]
  input  [31:0] io_in_B_1_12, // @[:@7775.4]
  input  [31:0] io_in_B_1_13, // @[:@7775.4]
  input  [31:0] io_in_B_1_14, // @[:@7775.4]
  input  [31:0] io_in_B_1_15, // @[:@7775.4]
  input  [31:0] io_in_B_2_0, // @[:@7775.4]
  input  [31:0] io_in_B_2_1, // @[:@7775.4]
  input  [31:0] io_in_B_2_2, // @[:@7775.4]
  input  [31:0] io_in_B_2_3, // @[:@7775.4]
  input  [31:0] io_in_B_2_4, // @[:@7775.4]
  input  [31:0] io_in_B_2_5, // @[:@7775.4]
  input  [31:0] io_in_B_2_6, // @[:@7775.4]
  input  [31:0] io_in_B_2_7, // @[:@7775.4]
  input  [31:0] io_in_B_2_8, // @[:@7775.4]
  input  [31:0] io_in_B_2_9, // @[:@7775.4]
  input  [31:0] io_in_B_2_10, // @[:@7775.4]
  input  [31:0] io_in_B_2_11, // @[:@7775.4]
  input  [31:0] io_in_B_2_12, // @[:@7775.4]
  input  [31:0] io_in_B_2_13, // @[:@7775.4]
  input  [31:0] io_in_B_2_14, // @[:@7775.4]
  input  [31:0] io_in_B_2_15, // @[:@7775.4]
  input  [31:0] io_in_B_3_0, // @[:@7775.4]
  input  [31:0] io_in_B_3_1, // @[:@7775.4]
  input  [31:0] io_in_B_3_2, // @[:@7775.4]
  input  [31:0] io_in_B_3_3, // @[:@7775.4]
  input  [31:0] io_in_B_3_4, // @[:@7775.4]
  input  [31:0] io_in_B_3_5, // @[:@7775.4]
  input  [31:0] io_in_B_3_6, // @[:@7775.4]
  input  [31:0] io_in_B_3_7, // @[:@7775.4]
  input  [31:0] io_in_B_3_8, // @[:@7775.4]
  input  [31:0] io_in_B_3_9, // @[:@7775.4]
  input  [31:0] io_in_B_3_10, // @[:@7775.4]
  input  [31:0] io_in_B_3_11, // @[:@7775.4]
  input  [31:0] io_in_B_3_12, // @[:@7775.4]
  input  [31:0] io_in_B_3_13, // @[:@7775.4]
  input  [31:0] io_in_B_3_14, // @[:@7775.4]
  input  [31:0] io_in_B_3_15, // @[:@7775.4]
  input  [31:0] io_in_B_4_0, // @[:@7775.4]
  input  [31:0] io_in_B_4_1, // @[:@7775.4]
  input  [31:0] io_in_B_4_2, // @[:@7775.4]
  input  [31:0] io_in_B_4_3, // @[:@7775.4]
  input  [31:0] io_in_B_4_4, // @[:@7775.4]
  input  [31:0] io_in_B_4_5, // @[:@7775.4]
  input  [31:0] io_in_B_4_6, // @[:@7775.4]
  input  [31:0] io_in_B_4_7, // @[:@7775.4]
  input  [31:0] io_in_B_4_8, // @[:@7775.4]
  input  [31:0] io_in_B_4_9, // @[:@7775.4]
  input  [31:0] io_in_B_4_10, // @[:@7775.4]
  input  [31:0] io_in_B_4_11, // @[:@7775.4]
  input  [31:0] io_in_B_4_12, // @[:@7775.4]
  input  [31:0] io_in_B_4_13, // @[:@7775.4]
  input  [31:0] io_in_B_4_14, // @[:@7775.4]
  input  [31:0] io_in_B_4_15, // @[:@7775.4]
  input  [31:0] io_in_B_5_0, // @[:@7775.4]
  input  [31:0] io_in_B_5_1, // @[:@7775.4]
  input  [31:0] io_in_B_5_2, // @[:@7775.4]
  input  [31:0] io_in_B_5_3, // @[:@7775.4]
  input  [31:0] io_in_B_5_4, // @[:@7775.4]
  input  [31:0] io_in_B_5_5, // @[:@7775.4]
  input  [31:0] io_in_B_5_6, // @[:@7775.4]
  input  [31:0] io_in_B_5_7, // @[:@7775.4]
  input  [31:0] io_in_B_5_8, // @[:@7775.4]
  input  [31:0] io_in_B_5_9, // @[:@7775.4]
  input  [31:0] io_in_B_5_10, // @[:@7775.4]
  input  [31:0] io_in_B_5_11, // @[:@7775.4]
  input  [31:0] io_in_B_5_12, // @[:@7775.4]
  input  [31:0] io_in_B_5_13, // @[:@7775.4]
  input  [31:0] io_in_B_5_14, // @[:@7775.4]
  input  [31:0] io_in_B_5_15, // @[:@7775.4]
  input  [31:0] io_in_B_6_0, // @[:@7775.4]
  input  [31:0] io_in_B_6_1, // @[:@7775.4]
  input  [31:0] io_in_B_6_2, // @[:@7775.4]
  input  [31:0] io_in_B_6_3, // @[:@7775.4]
  input  [31:0] io_in_B_6_4, // @[:@7775.4]
  input  [31:0] io_in_B_6_5, // @[:@7775.4]
  input  [31:0] io_in_B_6_6, // @[:@7775.4]
  input  [31:0] io_in_B_6_7, // @[:@7775.4]
  input  [31:0] io_in_B_6_8, // @[:@7775.4]
  input  [31:0] io_in_B_6_9, // @[:@7775.4]
  input  [31:0] io_in_B_6_10, // @[:@7775.4]
  input  [31:0] io_in_B_6_11, // @[:@7775.4]
  input  [31:0] io_in_B_6_12, // @[:@7775.4]
  input  [31:0] io_in_B_6_13, // @[:@7775.4]
  input  [31:0] io_in_B_6_14, // @[:@7775.4]
  input  [31:0] io_in_B_6_15, // @[:@7775.4]
  input  [31:0] io_in_B_7_0, // @[:@7775.4]
  input  [31:0] io_in_B_7_1, // @[:@7775.4]
  input  [31:0] io_in_B_7_2, // @[:@7775.4]
  input  [31:0] io_in_B_7_3, // @[:@7775.4]
  input  [31:0] io_in_B_7_4, // @[:@7775.4]
  input  [31:0] io_in_B_7_5, // @[:@7775.4]
  input  [31:0] io_in_B_7_6, // @[:@7775.4]
  input  [31:0] io_in_B_7_7, // @[:@7775.4]
  input  [31:0] io_in_B_7_8, // @[:@7775.4]
  input  [31:0] io_in_B_7_9, // @[:@7775.4]
  input  [31:0] io_in_B_7_10, // @[:@7775.4]
  input  [31:0] io_in_B_7_11, // @[:@7775.4]
  input  [31:0] io_in_B_7_12, // @[:@7775.4]
  input  [31:0] io_in_B_7_13, // @[:@7775.4]
  input  [31:0] io_in_B_7_14, // @[:@7775.4]
  input  [31:0] io_in_B_7_15, // @[:@7775.4]
  input         io_in_cal, // @[:@7775.4]
  output [31:0] io_out_C_0_0, // @[:@7775.4]
  output [31:0] io_out_C_0_1, // @[:@7775.4]
  output [31:0] io_out_C_0_2, // @[:@7775.4]
  output [31:0] io_out_C_0_3, // @[:@7775.4]
  output [31:0] io_out_C_0_4, // @[:@7775.4]
  output [31:0] io_out_C_0_5, // @[:@7775.4]
  output [31:0] io_out_C_0_6, // @[:@7775.4]
  output [31:0] io_out_C_0_7, // @[:@7775.4]
  output [31:0] io_out_C_1_0, // @[:@7775.4]
  output [31:0] io_out_C_1_1, // @[:@7775.4]
  output [31:0] io_out_C_1_2, // @[:@7775.4]
  output [31:0] io_out_C_1_3, // @[:@7775.4]
  output [31:0] io_out_C_1_4, // @[:@7775.4]
  output [31:0] io_out_C_1_5, // @[:@7775.4]
  output [31:0] io_out_C_1_6, // @[:@7775.4]
  output [31:0] io_out_C_1_7, // @[:@7775.4]
  output [31:0] io_out_C_2_0, // @[:@7775.4]
  output [31:0] io_out_C_2_1, // @[:@7775.4]
  output [31:0] io_out_C_2_2, // @[:@7775.4]
  output [31:0] io_out_C_2_3, // @[:@7775.4]
  output [31:0] io_out_C_2_4, // @[:@7775.4]
  output [31:0] io_out_C_2_5, // @[:@7775.4]
  output [31:0] io_out_C_2_6, // @[:@7775.4]
  output [31:0] io_out_C_2_7, // @[:@7775.4]
  output [31:0] io_out_C_3_0, // @[:@7775.4]
  output [31:0] io_out_C_3_1, // @[:@7775.4]
  output [31:0] io_out_C_3_2, // @[:@7775.4]
  output [31:0] io_out_C_3_3, // @[:@7775.4]
  output [31:0] io_out_C_3_4, // @[:@7775.4]
  output [31:0] io_out_C_3_5, // @[:@7775.4]
  output [31:0] io_out_C_3_6, // @[:@7775.4]
  output [31:0] io_out_C_3_7, // @[:@7775.4]
  output        io_out_cal // @[:@7775.4]
);
  wire  TPU_clock; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_reset; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_A_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_2_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_in_B_3_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_2_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_tag_3_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_in_cal; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_A_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_2_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_B_3_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_0_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_1_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_2_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_4; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_5; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_6; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_tag_3_7; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_0_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_0_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_0_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_0_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_1_0; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_1_1; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_1_2; // @[STA_VDBB.scala 97:36:@8674.4]
  wire [31:0] TPU_io_out_result_1_3; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_io_out_cal; // @[STA_VDBB.scala 97:36:@8674.4]
  wire  TPU_1_clock; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_reset; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_A_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_2_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_in_B_3_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_2_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_tag_3_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_in_cal; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_A_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_2_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_B_3_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_0_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_1_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_2_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_4; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_5; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_6; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_tag_3_7; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_0_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_0_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_0_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_0_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_1_0; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_1_1; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_1_2; // @[STA_VDBB.scala 97:36:@8677.4]
  wire [31:0] TPU_1_io_out_result_1_3; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_1_io_out_cal; // @[STA_VDBB.scala 97:36:@8677.4]
  wire  TPU_2_clock; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_reset; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_A_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_2_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_in_B_3_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_2_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_tag_3_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_in_cal; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_A_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_2_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_B_3_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_0_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_1_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_2_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_4; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_5; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_6; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_tag_3_7; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_0_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_0_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_0_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_0_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_1_0; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_1_1; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_1_2; // @[STA_VDBB.scala 97:36:@8680.4]
  wire [31:0] TPU_2_io_out_result_1_3; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_2_io_out_cal; // @[STA_VDBB.scala 97:36:@8680.4]
  wire  TPU_3_clock; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_reset; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_A_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_2_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_in_B_3_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_2_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_tag_3_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_in_cal; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_A_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_2_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_B_3_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_0_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_1_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_2_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_4; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_5; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_6; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_tag_3_7; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_0_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_0_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_0_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_0_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_1_0; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_1_1; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_1_2; // @[STA_VDBB.scala 97:36:@8683.4]
  wire [31:0] TPU_3_io_out_result_1_3; // @[STA_VDBB.scala 97:36:@8683.4]
  wire  TPU_3_io_out_cal; // @[STA_VDBB.scala 97:36:@8683.4]
  reg [31:0] reg_A_1_0_0; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_0;
  reg [31:0] reg_A_1_0_1; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_1;
  reg [31:0] reg_A_1_0_2; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_2;
  reg [31:0] reg_A_1_0_3; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_3;
  reg [31:0] reg_A_1_0_4; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_4;
  reg [31:0] reg_A_1_0_5; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_5;
  reg [31:0] reg_A_1_0_6; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_6;
  reg [31:0] reg_A_1_0_7; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_7;
  reg [31:0] reg_A_1_1_0; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_8;
  reg [31:0] reg_A_1_1_1; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_9;
  reg [31:0] reg_A_1_1_2; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_10;
  reg [31:0] reg_A_1_1_3; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_11;
  reg [31:0] reg_A_1_1_4; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_12;
  reg [31:0] reg_A_1_1_5; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_13;
  reg [31:0] reg_A_1_1_6; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_14;
  reg [31:0] reg_A_1_1_7; // @[STA_VDBB.scala 61:24:@7812.4]
  reg [31:0] _RAND_15;
  reg [31:0] reg_A_2_0_0; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_16;
  reg [31:0] reg_A_2_0_1; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_17;
  reg [31:0] reg_A_2_0_2; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_18;
  reg [31:0] reg_A_2_0_3; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_19;
  reg [31:0] reg_A_2_0_4; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_20;
  reg [31:0] reg_A_2_0_5; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_21;
  reg [31:0] reg_A_2_0_6; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_22;
  reg [31:0] reg_A_2_0_7; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_23;
  reg [31:0] reg_A_2_1_0; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_24;
  reg [31:0] reg_A_2_1_1; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_25;
  reg [31:0] reg_A_2_1_2; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_26;
  reg [31:0] reg_A_2_1_3; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_27;
  reg [31:0] reg_A_2_1_4; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_28;
  reg [31:0] reg_A_2_1_5; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_29;
  reg [31:0] reg_A_2_1_6; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_30;
  reg [31:0] reg_A_2_1_7; // @[STA_VDBB.scala 62:24:@7848.4]
  reg [31:0] _RAND_31;
  reg [31:0] reg_A_3_0_0; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_32;
  reg [31:0] reg_A_3_0_1; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_33;
  reg [31:0] reg_A_3_0_2; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_34;
  reg [31:0] reg_A_3_0_3; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_35;
  reg [31:0] reg_A_3_0_4; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_36;
  reg [31:0] reg_A_3_0_5; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_37;
  reg [31:0] reg_A_3_0_6; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_38;
  reg [31:0] reg_A_3_0_7; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_39;
  reg [31:0] reg_A_3_1_0; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_40;
  reg [31:0] reg_A_3_1_1; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_41;
  reg [31:0] reg_A_3_1_2; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_42;
  reg [31:0] reg_A_3_1_3; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_43;
  reg [31:0] reg_A_3_1_4; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_44;
  reg [31:0] reg_A_3_1_5; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_45;
  reg [31:0] reg_A_3_1_6; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_46;
  reg [31:0] reg_A_3_1_7; // @[STA_VDBB.scala 63:24:@7884.4]
  reg [31:0] _RAND_47;
  reg [31:0] reg_A_4_0_0; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_48;
  reg [31:0] reg_A_4_0_1; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_49;
  reg [31:0] reg_A_4_0_2; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_50;
  reg [31:0] reg_A_4_0_3; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_51;
  reg [31:0] reg_A_4_0_4; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_52;
  reg [31:0] reg_A_4_0_5; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_53;
  reg [31:0] reg_A_4_0_6; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_54;
  reg [31:0] reg_A_4_0_7; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_55;
  reg [31:0] reg_A_4_1_0; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_56;
  reg [31:0] reg_A_4_1_1; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_57;
  reg [31:0] reg_A_4_1_2; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_58;
  reg [31:0] reg_A_4_1_3; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_59;
  reg [31:0] reg_A_4_1_4; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_60;
  reg [31:0] reg_A_4_1_5; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_61;
  reg [31:0] reg_A_4_1_6; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_62;
  reg [31:0] reg_A_4_1_7; // @[STA_VDBB.scala 64:24:@7920.4]
  reg [31:0] _RAND_63;
  reg [31:0] reg_B_1_0_0; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_64;
  reg [31:0] reg_B_1_0_1; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_65;
  reg [31:0] reg_B_1_0_2; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_66;
  reg [31:0] reg_B_1_0_3; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_67;
  reg [31:0] reg_B_1_0_4; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_68;
  reg [31:0] reg_B_1_0_5; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_69;
  reg [31:0] reg_B_1_0_6; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_70;
  reg [31:0] reg_B_1_0_7; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_71;
  reg [31:0] reg_B_1_1_0; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_72;
  reg [31:0] reg_B_1_1_1; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_73;
  reg [31:0] reg_B_1_1_2; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_74;
  reg [31:0] reg_B_1_1_3; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_75;
  reg [31:0] reg_B_1_1_4; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_76;
  reg [31:0] reg_B_1_1_5; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_77;
  reg [31:0] reg_B_1_1_6; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_78;
  reg [31:0] reg_B_1_1_7; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_79;
  reg [31:0] reg_B_1_2_0; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_80;
  reg [31:0] reg_B_1_2_1; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_81;
  reg [31:0] reg_B_1_2_2; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_82;
  reg [31:0] reg_B_1_2_3; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_83;
  reg [31:0] reg_B_1_2_4; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_84;
  reg [31:0] reg_B_1_2_5; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_85;
  reg [31:0] reg_B_1_2_6; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_86;
  reg [31:0] reg_B_1_2_7; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_87;
  reg [31:0] reg_B_1_3_0; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_88;
  reg [31:0] reg_B_1_3_1; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_89;
  reg [31:0] reg_B_1_3_2; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_90;
  reg [31:0] reg_B_1_3_3; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_91;
  reg [31:0] reg_B_1_3_4; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_92;
  reg [31:0] reg_B_1_3_5; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_93;
  reg [31:0] reg_B_1_3_6; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_94;
  reg [31:0] reg_B_1_3_7; // @[STA_VDBB.scala 75:24:@8054.4]
  reg [31:0] _RAND_95;
  reg [31:0] reg_B_2_0_0; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_96;
  reg [31:0] reg_B_2_0_1; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_97;
  reg [31:0] reg_B_2_0_2; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_98;
  reg [31:0] reg_B_2_0_3; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_99;
  reg [31:0] reg_B_2_0_4; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_100;
  reg [31:0] reg_B_2_0_5; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_101;
  reg [31:0] reg_B_2_0_6; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_102;
  reg [31:0] reg_B_2_0_7; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_103;
  reg [31:0] reg_B_2_1_0; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_104;
  reg [31:0] reg_B_2_1_1; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_105;
  reg [31:0] reg_B_2_1_2; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_106;
  reg [31:0] reg_B_2_1_3; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_107;
  reg [31:0] reg_B_2_1_4; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_108;
  reg [31:0] reg_B_2_1_5; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_109;
  reg [31:0] reg_B_2_1_6; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_110;
  reg [31:0] reg_B_2_1_7; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_111;
  reg [31:0] reg_B_2_2_0; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_112;
  reg [31:0] reg_B_2_2_1; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_113;
  reg [31:0] reg_B_2_2_2; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_114;
  reg [31:0] reg_B_2_2_3; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_115;
  reg [31:0] reg_B_2_2_4; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_116;
  reg [31:0] reg_B_2_2_5; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_117;
  reg [31:0] reg_B_2_2_6; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_118;
  reg [31:0] reg_B_2_2_7; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_119;
  reg [31:0] reg_B_2_3_0; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_120;
  reg [31:0] reg_B_2_3_1; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_121;
  reg [31:0] reg_B_2_3_2; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_122;
  reg [31:0] reg_B_2_3_3; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_123;
  reg [31:0] reg_B_2_3_4; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_124;
  reg [31:0] reg_B_2_3_5; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_125;
  reg [31:0] reg_B_2_3_6; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_126;
  reg [31:0] reg_B_2_3_7; // @[STA_VDBB.scala 76:24:@8124.4]
  reg [31:0] _RAND_127;
  reg [31:0] reg_B_3_0_0; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_128;
  reg [31:0] reg_B_3_0_1; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_129;
  reg [31:0] reg_B_3_0_2; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_130;
  reg [31:0] reg_B_3_0_3; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_131;
  reg [31:0] reg_B_3_0_4; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_132;
  reg [31:0] reg_B_3_0_5; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_133;
  reg [31:0] reg_B_3_0_6; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_134;
  reg [31:0] reg_B_3_0_7; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_135;
  reg [31:0] reg_B_3_1_0; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_136;
  reg [31:0] reg_B_3_1_1; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_137;
  reg [31:0] reg_B_3_1_2; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_138;
  reg [31:0] reg_B_3_1_3; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_139;
  reg [31:0] reg_B_3_1_4; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_140;
  reg [31:0] reg_B_3_1_5; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_141;
  reg [31:0] reg_B_3_1_6; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_142;
  reg [31:0] reg_B_3_1_7; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_143;
  reg [31:0] reg_B_3_2_0; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_144;
  reg [31:0] reg_B_3_2_1; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_145;
  reg [31:0] reg_B_3_2_2; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_146;
  reg [31:0] reg_B_3_2_3; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_147;
  reg [31:0] reg_B_3_2_4; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_148;
  reg [31:0] reg_B_3_2_5; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_149;
  reg [31:0] reg_B_3_2_6; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_150;
  reg [31:0] reg_B_3_2_7; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_151;
  reg [31:0] reg_B_3_3_0; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_152;
  reg [31:0] reg_B_3_3_1; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_153;
  reg [31:0] reg_B_3_3_2; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_154;
  reg [31:0] reg_B_3_3_3; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_155;
  reg [31:0] reg_B_3_3_4; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_156;
  reg [31:0] reg_B_3_3_5; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_157;
  reg [31:0] reg_B_3_3_6; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_158;
  reg [31:0] reg_B_3_3_7; // @[STA_VDBB.scala 77:24:@8194.4]
  reg [31:0] _RAND_159;
  reg [31:0] reg_B_4_0_0; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_160;
  reg [31:0] reg_B_4_0_1; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_161;
  reg [31:0] reg_B_4_0_2; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_162;
  reg [31:0] reg_B_4_0_3; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_163;
  reg [31:0] reg_B_4_0_4; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_164;
  reg [31:0] reg_B_4_0_5; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_165;
  reg [31:0] reg_B_4_0_6; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_166;
  reg [31:0] reg_B_4_0_7; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_167;
  reg [31:0] reg_B_4_1_0; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_168;
  reg [31:0] reg_B_4_1_1; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_169;
  reg [31:0] reg_B_4_1_2; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_170;
  reg [31:0] reg_B_4_1_3; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_171;
  reg [31:0] reg_B_4_1_4; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_172;
  reg [31:0] reg_B_4_1_5; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_173;
  reg [31:0] reg_B_4_1_6; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_174;
  reg [31:0] reg_B_4_1_7; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_175;
  reg [31:0] reg_B_4_2_0; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_176;
  reg [31:0] reg_B_4_2_1; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_177;
  reg [31:0] reg_B_4_2_2; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_178;
  reg [31:0] reg_B_4_2_3; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_179;
  reg [31:0] reg_B_4_2_4; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_180;
  reg [31:0] reg_B_4_2_5; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_181;
  reg [31:0] reg_B_4_2_6; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_182;
  reg [31:0] reg_B_4_2_7; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_183;
  reg [31:0] reg_B_4_3_0; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_184;
  reg [31:0] reg_B_4_3_1; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_185;
  reg [31:0] reg_B_4_3_2; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_186;
  reg [31:0] reg_B_4_3_3; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_187;
  reg [31:0] reg_B_4_3_4; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_188;
  reg [31:0] reg_B_4_3_5; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_189;
  reg [31:0] reg_B_4_3_6; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_190;
  reg [31:0] reg_B_4_3_7; // @[STA_VDBB.scala 78:24:@8264.4]
  reg [31:0] _RAND_191;
  reg  cal_state_0; // @[STA_VDBB.scala 113:26:@9855.4]
  reg [31:0] _RAND_192;
  reg  cal_state_1; // @[STA_VDBB.scala 113:26:@9855.4]
  reg [31:0] _RAND_193;
  reg  cal_state_2; // @[STA_VDBB.scala 113:26:@9855.4]
  reg [31:0] _RAND_194;
  wire  TPUs_1_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8857.4]
  wire  TPUs_2_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9027.4]
  wire  _T_40965; // @[STA_VDBB.scala 115:35:@9857.4]
  wire  _T_40966; // @[STA_VDBB.scala 117:30:@9860.4]
  reg [31:0] result_0_0; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_195;
  reg [31:0] result_0_1; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_196;
  reg [31:0] result_0_2; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_197;
  reg [31:0] result_0_3; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_198;
  reg [31:0] result_0_4; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_199;
  reg [31:0] result_0_5; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_200;
  reg [31:0] result_0_6; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_201;
  reg [31:0] result_0_7; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_202;
  reg [31:0] result_1_0; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_203;
  reg [31:0] result_1_1; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_204;
  reg [31:0] result_1_2; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_205;
  reg [31:0] result_1_3; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_206;
  reg [31:0] result_1_4; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_207;
  reg [31:0] result_1_5; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_208;
  reg [31:0] result_1_6; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_209;
  reg [31:0] result_1_7; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_210;
  reg [31:0] result_2_0; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_211;
  reg [31:0] result_2_1; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_212;
  reg [31:0] result_2_2; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_213;
  reg [31:0] result_2_3; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_214;
  reg [31:0] result_2_4; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_215;
  reg [31:0] result_2_5; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_216;
  reg [31:0] result_2_6; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_217;
  reg [31:0] result_2_7; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_218;
  reg [31:0] result_3_0; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_219;
  reg [31:0] result_3_1; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_220;
  reg [31:0] result_3_2; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_221;
  reg [31:0] result_3_3; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_222;
  reg [31:0] result_3_4; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_223;
  reg [31:0] result_3_5; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_224;
  reg [31:0] result_3_6; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_225;
  reg [31:0] result_3_7; // @[STA_VDBB.scala 119:23:@9932.4]
  reg [31:0] _RAND_226;
  reg  cal_control_0; // @[STA_VDBB.scala 130:28:@10001.4]
  reg [31:0] _RAND_227;
  reg  cal_control_1; // @[STA_VDBB.scala 130:28:@10001.4]
  reg [31:0] _RAND_228;
  reg  cal_control_2; // @[STA_VDBB.scala 130:28:@10001.4]
  reg [31:0] _RAND_229;
  reg [2:0] stateReg; // @[STA_VDBB.scala 138:25:@10006.4]
  reg [31:0] _RAND_230;
  reg  loop_reg; // @[STA_VDBB.scala 139:25:@10007.4]
  reg [31:0] _RAND_231;
  wire  _T_43000; // @[Conditional.scala 37:30:@10008.4]
  reg  _T_43002; // @[STA_VDBB.scala 143:32:@10010.6]
  reg [31:0] _RAND_232;
  wire  _T_43004; // @[STA_VDBB.scala 143:24:@10012.6]
  wire  _T_43005; // @[STA_VDBB.scala 143:22:@10013.6]
  wire [2:0] _GEN_0; // @[STA_VDBB.scala 143:44:@10014.6]
  wire  _T_43006; // @[Conditional.scala 37:30:@10019.6]
  wire  _T_43007; // @[Conditional.scala 37:30:@10021.8]
  wire  _GEN_1; // @[STA_VDBB.scala 159:29:@10141.12]
  wire [2:0] _GEN_2; // @[STA_VDBB.scala 159:29:@10141.12]
  wire  _GEN_3; // @[STA_VDBB.scala 159:29:@10141.12]
  wire  _GEN_4; // @[Conditional.scala 39:67:@10139.10]
  wire [2:0] _GEN_5; // @[Conditional.scala 39:67:@10139.10]
  wire  _GEN_6; // @[Conditional.scala 39:67:@10139.10]
  wire [31:0] _GEN_7; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_8; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_9; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_10; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_11; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_12; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_13; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_14; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_15; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_16; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_17; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_18; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_19; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_20; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_21; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_22; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_23; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_24; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_25; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_26; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_27; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_28; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_29; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_30; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_31; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_32; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_33; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_34; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_35; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_36; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_37; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_38; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_39; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_40; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_41; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_42; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_43; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_44; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_45; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_46; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_47; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_48; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_49; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_50; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_51; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_52; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_53; // @[Conditional.scala 40:58:@10022.8]
  wire [31:0] _GEN_54; // @[Conditional.scala 40:58:@10022.8]
  wire  _GEN_119; // @[Conditional.scala 40:58:@10022.8]
  wire  _GEN_120; // @[Conditional.scala 40:58:@10022.8]
  wire [2:0] _GEN_121; // @[Conditional.scala 40:58:@10022.8]
  wire  _T_43011; // @[Conditional.scala 37:30:@10149.8]
  wire  _GEN_122; // @[STA_VDBB.scala 179:29:@10271.14]
  wire [2:0] _GEN_123; // @[STA_VDBB.scala 179:29:@10271.14]
  wire  _GEN_124; // @[STA_VDBB.scala 179:29:@10271.14]
  wire  _GEN_125; // @[Conditional.scala 39:67:@10269.12]
  wire [2:0] _GEN_126; // @[Conditional.scala 39:67:@10269.12]
  wire  _GEN_127; // @[Conditional.scala 39:67:@10269.12]
  wire [31:0] TPUs_0_out_A_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8760.4]
  wire [31:0] _GEN_128; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8761.4]
  wire [31:0] _GEN_129; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8762.4]
  wire [31:0] _GEN_130; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8763.4]
  wire [31:0] _GEN_131; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8764.4]
  wire [31:0] _GEN_132; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8765.4]
  wire [31:0] _GEN_133; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8766.4]
  wire [31:0] _GEN_134; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8767.4]
  wire [31:0] _GEN_135; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8768.4]
  wire [31:0] _GEN_136; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8769.4]
  wire [31:0] _GEN_137; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8770.4]
  wire [31:0] _GEN_138; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8771.4]
  wire [31:0] _GEN_139; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8772.4]
  wire [31:0] _GEN_140; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8773.4]
  wire [31:0] _GEN_141; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8774.4]
  wire [31:0] _GEN_142; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_A_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8775.4]
  wire [31:0] _GEN_143; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8728.4]
  wire [31:0] _GEN_144; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8729.4]
  wire [31:0] _GEN_145; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8730.4]
  wire [31:0] _GEN_146; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8731.4]
  wire [31:0] _GEN_147; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8732.4]
  wire [31:0] _GEN_148; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8733.4]
  wire [31:0] _GEN_149; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8734.4]
  wire [31:0] _GEN_150; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8735.4]
  wire [31:0] _GEN_151; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8736.4]
  wire [31:0] _GEN_152; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8737.4]
  wire [31:0] _GEN_153; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8738.4]
  wire [31:0] _GEN_154; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8739.4]
  wire [31:0] _GEN_155; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8740.4]
  wire [31:0] _GEN_156; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8741.4]
  wire [31:0] _GEN_157; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8742.4]
  wire [31:0] _GEN_158; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8743.4]
  wire [31:0] _GEN_159; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8744.4]
  wire [31:0] _GEN_160; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8745.4]
  wire [31:0] _GEN_161; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8746.4]
  wire [31:0] _GEN_162; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8747.4]
  wire [31:0] _GEN_163; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8748.4]
  wire [31:0] _GEN_164; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8749.4]
  wire [31:0] _GEN_165; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8750.4]
  wire [31:0] _GEN_166; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_2_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8751.4]
  wire [31:0] _GEN_167; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8752.4]
  wire [31:0] _GEN_168; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8753.4]
  wire [31:0] _GEN_169; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8754.4]
  wire [31:0] _GEN_170; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8755.4]
  wire [31:0] _GEN_171; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8756.4]
  wire [31:0] _GEN_172; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8757.4]
  wire [31:0] _GEN_173; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8758.4]
  wire [31:0] _GEN_174; // @[Conditional.scala 40:58:@10152.10]
  wire [31:0] TPUs_0_out_B_3_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8759.4]
  wire [31:0] _GEN_175; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8696.4]
  wire  _GEN_208; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8697.4]
  wire  _GEN_209; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8698.4]
  wire  _GEN_210; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8699.4]
  wire  _GEN_211; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8700.4]
  wire  _GEN_212; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8701.4]
  wire  _GEN_213; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8702.4]
  wire  _GEN_214; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8703.4]
  wire  _GEN_215; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8704.4]
  wire  _GEN_216; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8705.4]
  wire  _GEN_217; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8706.4]
  wire  _GEN_218; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8707.4]
  wire  _GEN_219; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8708.4]
  wire  _GEN_220; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8709.4]
  wire  _GEN_221; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8710.4]
  wire  _GEN_222; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8711.4]
  wire  _GEN_223; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8712.4]
  wire  _GEN_224; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8713.4]
  wire  _GEN_225; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8714.4]
  wire  _GEN_226; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8715.4]
  wire  _GEN_227; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8716.4]
  wire  _GEN_228; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8717.4]
  wire  _GEN_229; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8718.4]
  wire  _GEN_230; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_2_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8719.4]
  wire  _GEN_231; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8720.4]
  wire  _GEN_232; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8721.4]
  wire  _GEN_233; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8722.4]
  wire  _GEN_234; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8723.4]
  wire  _GEN_235; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8724.4]
  wire  _GEN_236; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8725.4]
  wire  _GEN_237; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8726.4]
  wire  _GEN_238; // @[Conditional.scala 40:58:@10152.10]
  wire  TPUs_0_out_tag_3_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8727.4]
  wire  _GEN_239; // @[Conditional.scala 40:58:@10152.10]
  wire  _GEN_240; // @[Conditional.scala 40:58:@10152.10]
  wire  _GEN_241; // @[Conditional.scala 40:58:@10152.10]
  wire [2:0] _GEN_242; // @[Conditional.scala 40:58:@10152.10]
  wire  _T_43016; // @[Conditional.scala 37:30:@10279.10]
  wire  _T_43021; // @[STA_VDBB.scala 200:29:@10402.16]
  wire  _GEN_243; // @[STA_VDBB.scala 200:45:@10403.16]
  wire [2:0] _GEN_244; // @[STA_VDBB.scala 200:45:@10403.16]
  wire  _GEN_245; // @[STA_VDBB.scala 200:45:@10403.16]
  wire  _GEN_246; // @[Conditional.scala 39:67:@10399.14]
  wire  _GEN_247; // @[Conditional.scala 39:67:@10399.14]
  wire [2:0] _GEN_248; // @[Conditional.scala 39:67:@10399.14]
  wire  _GEN_249; // @[Conditional.scala 39:67:@10399.14]
  wire [31:0] _GEN_250; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_251; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_252; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_253; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_254; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_255; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_256; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_257; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_258; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_259; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_260; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_261; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_262; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_263; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_264; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_265; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_266; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_267; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_268; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_269; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_270; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_271; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_272; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_273; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_274; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_275; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_276; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_277; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_278; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_279; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_280; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_281; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_282; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_283; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_284; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_285; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_286; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_287; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_288; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_289; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_290; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_291; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_292; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_293; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_294; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_295; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_296; // @[Conditional.scala 40:58:@10282.12]
  wire [31:0] _GEN_297; // @[Conditional.scala 40:58:@10282.12]
  wire  _GEN_362; // @[Conditional.scala 40:58:@10282.12]
  wire  _GEN_363; // @[Conditional.scala 40:58:@10282.12]
  wire  _GEN_364; // @[Conditional.scala 40:58:@10282.12]
  wire [2:0] _GEN_365; // @[Conditional.scala 40:58:@10282.12]
  wire  _T_43024; // @[Conditional.scala 37:30:@10412.12]
  wire [2:0] _GEN_366; // @[STA_VDBB.scala 221:29:@10534.18]
  wire [2:0] _GEN_368; // @[Conditional.scala 39:67:@10532.16]
  wire [31:0] _GEN_370; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_371; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_372; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_373; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_374; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_375; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_376; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_377; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_378; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_379; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_380; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_381; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_382; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_383; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_384; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_385; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_386; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_387; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_388; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_389; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_390; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_391; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_392; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_393; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_394; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_395; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_396; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_397; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_398; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_399; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_400; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_401; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_402; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_403; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_404; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_405; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_406; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_407; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_408; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_409; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_410; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_411; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_412; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_413; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_414; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_415; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_416; // @[Conditional.scala 40:58:@10415.14]
  wire [31:0] _GEN_417; // @[Conditional.scala 40:58:@10415.14]
  wire [2:0] _GEN_484; // @[Conditional.scala 40:58:@10415.14]
  wire  _T_43029; // @[Conditional.scala 37:30:@10542.14]
  wire  _GEN_485; // @[STA_VDBB.scala 237:29:@10552.20]
  wire [2:0] _GEN_486; // @[STA_VDBB.scala 237:29:@10552.20]
  wire  _GEN_487; // @[STA_VDBB.scala 237:29:@10552.20]
  wire  _GEN_488; // @[Conditional.scala 39:67:@10550.18]
  wire  _GEN_489; // @[Conditional.scala 39:67:@10550.18]
  wire [2:0] _GEN_490; // @[Conditional.scala 39:67:@10550.18]
  wire  _GEN_491; // @[Conditional.scala 39:67:@10550.18]
  wire  _GEN_492; // @[Conditional.scala 40:58:@10545.16]
  wire  _GEN_493; // @[Conditional.scala 40:58:@10545.16]
  wire  _GEN_494; // @[Conditional.scala 40:58:@10545.16]
  wire [2:0] _GEN_495; // @[Conditional.scala 40:58:@10545.16]
  wire  _GEN_496; // @[Conditional.scala 39:67:@10543.14]
  wire  _GEN_497; // @[Conditional.scala 39:67:@10543.14]
  wire  _GEN_498; // @[Conditional.scala 39:67:@10543.14]
  wire [2:0] _GEN_499; // @[Conditional.scala 39:67:@10543.14]
  wire [31:0] _GEN_500; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_501; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_502; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_503; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_504; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_505; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_506; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_507; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_508; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_509; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_510; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_511; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_512; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_513; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_514; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_515; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_516; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_517; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_518; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_519; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_520; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_521; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_522; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_523; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_524; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_525; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_526; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_527; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_528; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_529; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_530; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_531; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_532; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_533; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_534; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_535; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_536; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_537; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_538; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_539; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_540; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_541; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_542; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_543; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_544; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_545; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_546; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_547; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_580; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_581; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_582; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_583; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_584; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_585; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_586; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_587; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_588; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_589; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_590; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_591; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_592; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_593; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_594; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_595; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_596; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_597; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_598; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_599; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_600; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_601; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_602; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_603; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_604; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_605; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_606; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_607; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_608; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_609; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_610; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_611; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_612; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_613; // @[Conditional.scala 39:67:@10413.12]
  wire [2:0] _GEN_614; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_615; // @[Conditional.scala 39:67:@10413.12]
  wire  _GEN_616; // @[Conditional.scala 39:67:@10413.12]
  wire [31:0] _GEN_617; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_618; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_619; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_620; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_621; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_622; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_623; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_624; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_625; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_626; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_627; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_628; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_629; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_630; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_631; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_632; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_633; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_634; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_635; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_636; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_637; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_638; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_639; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_640; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_641; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_642; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_643; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_644; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_645; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_646; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_647; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_648; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_649; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_650; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_651; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_652; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_653; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_654; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_655; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_656; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_657; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_658; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_659; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_660; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_661; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_662; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_663; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_664; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_729; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_730; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_731; // @[Conditional.scala 39:67:@10280.10]
  wire [2:0] _GEN_732; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_733; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_734; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_735; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_736; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_737; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_738; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_739; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_740; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_741; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_742; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_743; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_744; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_745; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_746; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_747; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_748; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_749; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_750; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_751; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_752; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_753; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_754; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_755; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_756; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_757; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_758; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_759; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_760; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_761; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_762; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_763; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_764; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_765; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_766; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_767; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_768; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_769; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_770; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_771; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_772; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_773; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_774; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_775; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_776; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_777; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_778; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_779; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_780; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_781; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_782; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_783; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_784; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_785; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_786; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_787; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_788; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_789; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_790; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_791; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_792; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_793; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_794; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_795; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_796; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_797; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_798; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_799; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_800; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_801; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_802; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_803; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_804; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_805; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_806; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_807; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_808; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_809; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_810; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_811; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_812; // @[Conditional.scala 39:67:@10280.10]
  wire  _GEN_813; // @[Conditional.scala 39:67:@10280.10]
  wire [31:0] _GEN_814; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_815; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_816; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_817; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_818; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_819; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_820; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_821; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_822; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_823; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_824; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_825; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_826; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_827; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_828; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_829; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_830; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_831; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_832; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_833; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_834; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_835; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_836; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_837; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_838; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_839; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_840; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_841; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_842; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_843; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_844; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_845; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_846; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_847; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_848; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_849; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_850; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_851; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_852; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_853; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_854; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_855; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_856; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_857; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_858; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_859; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_860; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_861; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_894; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_895; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_896; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_897; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_898; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_899; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_900; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_901; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_902; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_903; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_904; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_905; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_906; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_907; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_908; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_909; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_910; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_911; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_912; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_913; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_914; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_915; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_916; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_917; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_918; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_919; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_920; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_921; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_922; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_923; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_924; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_925; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_926; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_927; // @[Conditional.scala 39:67:@10150.8]
  wire [2:0] _GEN_928; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_929; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_930; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_931; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_932; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_933; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_934; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_935; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_936; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_937; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_938; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_939; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_940; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_941; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_942; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_943; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_944; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_945; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_946; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_947; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_948; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_949; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_950; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_951; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_952; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_953; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_954; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_955; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_956; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_957; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_958; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_959; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_960; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_961; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_962; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_963; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_964; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_965; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_966; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_967; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_968; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_969; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_970; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_971; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_972; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_973; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_974; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_975; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_976; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_1009; // @[Conditional.scala 39:67:@10150.8]
  wire  _GEN_1010; // @[Conditional.scala 39:67:@10150.8]
  wire [31:0] _GEN_1011; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1012; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1013; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1014; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1015; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1016; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1017; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1018; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1019; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1020; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1021; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1022; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1023; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1024; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1025; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1026; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1027; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1028; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1029; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1030; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1031; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1032; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1033; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1034; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1035; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1036; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1037; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1038; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1039; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1040; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1041; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1042; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1043; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1044; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1045; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1046; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1047; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1048; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1049; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1050; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1051; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1052; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1053; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1054; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1055; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1056; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1057; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1058; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1123; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1124; // @[Conditional.scala 39:67:@10020.6]
  wire [2:0] _GEN_1125; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1126; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1127; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1128; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1129; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1130; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1131; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1132; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1133; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1134; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1135; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1136; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1137; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1138; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1139; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1140; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1141; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1142; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1143; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1144; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1145; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1146; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1147; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1148; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1149; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1150; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1151; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1152; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1153; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1154; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1155; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1156; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1157; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1158; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1159; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1160; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1161; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1162; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1163; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1164; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1165; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1166; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1167; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1168; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1169; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1170; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1171; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1172; // @[Conditional.scala 39:67:@10020.6]
  wire [31:0] _GEN_1173; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1174; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1175; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1176; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1177; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1178; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1179; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1180; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1181; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1182; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1183; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1184; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1185; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1186; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1187; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1188; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1189; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1190; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1191; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1192; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1193; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1194; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1195; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1196; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1197; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1198; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1199; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1200; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1201; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1202; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1203; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1204; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1205; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1206; // @[Conditional.scala 39:67:@10020.6]
  wire  _GEN_1207; // @[Conditional.scala 39:67:@10020.6]
  wire [2:0] _GEN_1208; // @[Conditional.scala 40:58:@10009.4]
  wire  _GEN_1321; // @[Conditional.scala 40:58:@10009.4]
  wire  _GEN_1322; // @[Conditional.scala 40:58:@10009.4]
  wire  _GEN_1403; // @[Conditional.scala 40:58:@10009.4]
  wire  _GEN_1404; // @[Conditional.scala 40:58:@10009.4]
  wire [31:0] TPUs_0_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8688.4]
  wire [31:0] TPUs_0_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8689.4]
  wire [31:0] TPUs_0_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8690.4]
  wire [31:0] TPUs_0_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8691.4]
  wire [31:0] TPUs_0_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8692.4]
  wire [31:0] TPUs_0_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8693.4]
  wire [31:0] TPUs_0_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8694.4]
  wire [31:0] TPUs_0_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8695.4]
  wire  TPUs_0_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8687.4]
  wire [31:0] TPUs_1_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8858.4]
  wire [31:0] TPUs_1_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8859.4]
  wire [31:0] TPUs_1_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8860.4]
  wire [31:0] TPUs_1_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8861.4]
  wire [31:0] TPUs_1_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8862.4]
  wire [31:0] TPUs_1_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8863.4]
  wire [31:0] TPUs_1_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8864.4]
  wire [31:0] TPUs_1_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8865.4]
  wire [31:0] TPUs_2_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9028.4]
  wire [31:0] TPUs_2_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9029.4]
  wire [31:0] TPUs_2_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9030.4]
  wire [31:0] TPUs_2_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9031.4]
  wire [31:0] TPUs_2_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9032.4]
  wire [31:0] TPUs_2_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9033.4]
  wire [31:0] TPUs_2_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9034.4]
  wire [31:0] TPUs_2_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9035.4]
  wire [31:0] TPUs_3_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9198.4]
  wire [31:0] TPUs_3_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9199.4]
  wire [31:0] TPUs_3_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9200.4]
  wire [31:0] TPUs_3_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9201.4]
  wire [31:0] TPUs_3_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9202.4]
  wire [31:0] TPUs_3_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9203.4]
  wire [31:0] TPUs_3_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9204.4]
  wire [31:0] TPUs_3_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9205.4]
  wire  TPUs_3_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9197.4]
  TPU TPU ( // @[STA_VDBB.scala 97:36:@8674.4]
    .clock(TPU_clock),
    .reset(TPU_reset),
    .io_in_A_0_0(TPU_io_in_A_0_0),
    .io_in_A_0_1(TPU_io_in_A_0_1),
    .io_in_A_0_2(TPU_io_in_A_0_2),
    .io_in_A_0_3(TPU_io_in_A_0_3),
    .io_in_A_0_4(TPU_io_in_A_0_4),
    .io_in_A_0_5(TPU_io_in_A_0_5),
    .io_in_A_0_6(TPU_io_in_A_0_6),
    .io_in_A_0_7(TPU_io_in_A_0_7),
    .io_in_A_1_0(TPU_io_in_A_1_0),
    .io_in_A_1_1(TPU_io_in_A_1_1),
    .io_in_A_1_2(TPU_io_in_A_1_2),
    .io_in_A_1_3(TPU_io_in_A_1_3),
    .io_in_A_1_4(TPU_io_in_A_1_4),
    .io_in_A_1_5(TPU_io_in_A_1_5),
    .io_in_A_1_6(TPU_io_in_A_1_6),
    .io_in_A_1_7(TPU_io_in_A_1_7),
    .io_in_B_0_0(TPU_io_in_B_0_0),
    .io_in_B_0_1(TPU_io_in_B_0_1),
    .io_in_B_0_2(TPU_io_in_B_0_2),
    .io_in_B_0_3(TPU_io_in_B_0_3),
    .io_in_B_0_4(TPU_io_in_B_0_4),
    .io_in_B_0_5(TPU_io_in_B_0_5),
    .io_in_B_0_6(TPU_io_in_B_0_6),
    .io_in_B_0_7(TPU_io_in_B_0_7),
    .io_in_B_1_0(TPU_io_in_B_1_0),
    .io_in_B_1_1(TPU_io_in_B_1_1),
    .io_in_B_1_2(TPU_io_in_B_1_2),
    .io_in_B_1_3(TPU_io_in_B_1_3),
    .io_in_B_1_4(TPU_io_in_B_1_4),
    .io_in_B_1_5(TPU_io_in_B_1_5),
    .io_in_B_1_6(TPU_io_in_B_1_6),
    .io_in_B_1_7(TPU_io_in_B_1_7),
    .io_in_B_2_0(TPU_io_in_B_2_0),
    .io_in_B_2_1(TPU_io_in_B_2_1),
    .io_in_B_2_2(TPU_io_in_B_2_2),
    .io_in_B_2_3(TPU_io_in_B_2_3),
    .io_in_B_2_4(TPU_io_in_B_2_4),
    .io_in_B_2_5(TPU_io_in_B_2_5),
    .io_in_B_2_6(TPU_io_in_B_2_6),
    .io_in_B_2_7(TPU_io_in_B_2_7),
    .io_in_B_3_0(TPU_io_in_B_3_0),
    .io_in_B_3_1(TPU_io_in_B_3_1),
    .io_in_B_3_2(TPU_io_in_B_3_2),
    .io_in_B_3_3(TPU_io_in_B_3_3),
    .io_in_B_3_4(TPU_io_in_B_3_4),
    .io_in_B_3_5(TPU_io_in_B_3_5),
    .io_in_B_3_6(TPU_io_in_B_3_6),
    .io_in_B_3_7(TPU_io_in_B_3_7),
    .io_in_tag_0_0(TPU_io_in_tag_0_0),
    .io_in_tag_0_1(TPU_io_in_tag_0_1),
    .io_in_tag_0_2(TPU_io_in_tag_0_2),
    .io_in_tag_0_3(TPU_io_in_tag_0_3),
    .io_in_tag_0_4(TPU_io_in_tag_0_4),
    .io_in_tag_0_5(TPU_io_in_tag_0_5),
    .io_in_tag_0_6(TPU_io_in_tag_0_6),
    .io_in_tag_0_7(TPU_io_in_tag_0_7),
    .io_in_tag_1_0(TPU_io_in_tag_1_0),
    .io_in_tag_1_1(TPU_io_in_tag_1_1),
    .io_in_tag_1_2(TPU_io_in_tag_1_2),
    .io_in_tag_1_3(TPU_io_in_tag_1_3),
    .io_in_tag_1_4(TPU_io_in_tag_1_4),
    .io_in_tag_1_5(TPU_io_in_tag_1_5),
    .io_in_tag_1_6(TPU_io_in_tag_1_6),
    .io_in_tag_1_7(TPU_io_in_tag_1_7),
    .io_in_tag_2_0(TPU_io_in_tag_2_0),
    .io_in_tag_2_1(TPU_io_in_tag_2_1),
    .io_in_tag_2_2(TPU_io_in_tag_2_2),
    .io_in_tag_2_3(TPU_io_in_tag_2_3),
    .io_in_tag_2_4(TPU_io_in_tag_2_4),
    .io_in_tag_2_5(TPU_io_in_tag_2_5),
    .io_in_tag_2_6(TPU_io_in_tag_2_6),
    .io_in_tag_2_7(TPU_io_in_tag_2_7),
    .io_in_tag_3_0(TPU_io_in_tag_3_0),
    .io_in_tag_3_1(TPU_io_in_tag_3_1),
    .io_in_tag_3_2(TPU_io_in_tag_3_2),
    .io_in_tag_3_3(TPU_io_in_tag_3_3),
    .io_in_tag_3_4(TPU_io_in_tag_3_4),
    .io_in_tag_3_5(TPU_io_in_tag_3_5),
    .io_in_tag_3_6(TPU_io_in_tag_3_6),
    .io_in_tag_3_7(TPU_io_in_tag_3_7),
    .io_in_cal(TPU_io_in_cal),
    .io_out_A_0_0(TPU_io_out_A_0_0),
    .io_out_A_0_1(TPU_io_out_A_0_1),
    .io_out_A_0_2(TPU_io_out_A_0_2),
    .io_out_A_0_3(TPU_io_out_A_0_3),
    .io_out_A_0_4(TPU_io_out_A_0_4),
    .io_out_A_0_5(TPU_io_out_A_0_5),
    .io_out_A_0_6(TPU_io_out_A_0_6),
    .io_out_A_0_7(TPU_io_out_A_0_7),
    .io_out_A_1_0(TPU_io_out_A_1_0),
    .io_out_A_1_1(TPU_io_out_A_1_1),
    .io_out_A_1_2(TPU_io_out_A_1_2),
    .io_out_A_1_3(TPU_io_out_A_1_3),
    .io_out_A_1_4(TPU_io_out_A_1_4),
    .io_out_A_1_5(TPU_io_out_A_1_5),
    .io_out_A_1_6(TPU_io_out_A_1_6),
    .io_out_A_1_7(TPU_io_out_A_1_7),
    .io_out_B_0_0(TPU_io_out_B_0_0),
    .io_out_B_0_1(TPU_io_out_B_0_1),
    .io_out_B_0_2(TPU_io_out_B_0_2),
    .io_out_B_0_3(TPU_io_out_B_0_3),
    .io_out_B_0_4(TPU_io_out_B_0_4),
    .io_out_B_0_5(TPU_io_out_B_0_5),
    .io_out_B_0_6(TPU_io_out_B_0_6),
    .io_out_B_0_7(TPU_io_out_B_0_7),
    .io_out_B_1_0(TPU_io_out_B_1_0),
    .io_out_B_1_1(TPU_io_out_B_1_1),
    .io_out_B_1_2(TPU_io_out_B_1_2),
    .io_out_B_1_3(TPU_io_out_B_1_3),
    .io_out_B_1_4(TPU_io_out_B_1_4),
    .io_out_B_1_5(TPU_io_out_B_1_5),
    .io_out_B_1_6(TPU_io_out_B_1_6),
    .io_out_B_1_7(TPU_io_out_B_1_7),
    .io_out_B_2_0(TPU_io_out_B_2_0),
    .io_out_B_2_1(TPU_io_out_B_2_1),
    .io_out_B_2_2(TPU_io_out_B_2_2),
    .io_out_B_2_3(TPU_io_out_B_2_3),
    .io_out_B_2_4(TPU_io_out_B_2_4),
    .io_out_B_2_5(TPU_io_out_B_2_5),
    .io_out_B_2_6(TPU_io_out_B_2_6),
    .io_out_B_2_7(TPU_io_out_B_2_7),
    .io_out_B_3_0(TPU_io_out_B_3_0),
    .io_out_B_3_1(TPU_io_out_B_3_1),
    .io_out_B_3_2(TPU_io_out_B_3_2),
    .io_out_B_3_3(TPU_io_out_B_3_3),
    .io_out_B_3_4(TPU_io_out_B_3_4),
    .io_out_B_3_5(TPU_io_out_B_3_5),
    .io_out_B_3_6(TPU_io_out_B_3_6),
    .io_out_B_3_7(TPU_io_out_B_3_7),
    .io_out_tag_0_0(TPU_io_out_tag_0_0),
    .io_out_tag_0_1(TPU_io_out_tag_0_1),
    .io_out_tag_0_2(TPU_io_out_tag_0_2),
    .io_out_tag_0_3(TPU_io_out_tag_0_3),
    .io_out_tag_0_4(TPU_io_out_tag_0_4),
    .io_out_tag_0_5(TPU_io_out_tag_0_5),
    .io_out_tag_0_6(TPU_io_out_tag_0_6),
    .io_out_tag_0_7(TPU_io_out_tag_0_7),
    .io_out_tag_1_0(TPU_io_out_tag_1_0),
    .io_out_tag_1_1(TPU_io_out_tag_1_1),
    .io_out_tag_1_2(TPU_io_out_tag_1_2),
    .io_out_tag_1_3(TPU_io_out_tag_1_3),
    .io_out_tag_1_4(TPU_io_out_tag_1_4),
    .io_out_tag_1_5(TPU_io_out_tag_1_5),
    .io_out_tag_1_6(TPU_io_out_tag_1_6),
    .io_out_tag_1_7(TPU_io_out_tag_1_7),
    .io_out_tag_2_0(TPU_io_out_tag_2_0),
    .io_out_tag_2_1(TPU_io_out_tag_2_1),
    .io_out_tag_2_2(TPU_io_out_tag_2_2),
    .io_out_tag_2_3(TPU_io_out_tag_2_3),
    .io_out_tag_2_4(TPU_io_out_tag_2_4),
    .io_out_tag_2_5(TPU_io_out_tag_2_5),
    .io_out_tag_2_6(TPU_io_out_tag_2_6),
    .io_out_tag_2_7(TPU_io_out_tag_2_7),
    .io_out_tag_3_0(TPU_io_out_tag_3_0),
    .io_out_tag_3_1(TPU_io_out_tag_3_1),
    .io_out_tag_3_2(TPU_io_out_tag_3_2),
    .io_out_tag_3_3(TPU_io_out_tag_3_3),
    .io_out_tag_3_4(TPU_io_out_tag_3_4),
    .io_out_tag_3_5(TPU_io_out_tag_3_5),
    .io_out_tag_3_6(TPU_io_out_tag_3_6),
    .io_out_tag_3_7(TPU_io_out_tag_3_7),
    .io_out_result_0_0(TPU_io_out_result_0_0),
    .io_out_result_0_1(TPU_io_out_result_0_1),
    .io_out_result_0_2(TPU_io_out_result_0_2),
    .io_out_result_0_3(TPU_io_out_result_0_3),
    .io_out_result_1_0(TPU_io_out_result_1_0),
    .io_out_result_1_1(TPU_io_out_result_1_1),
    .io_out_result_1_2(TPU_io_out_result_1_2),
    .io_out_result_1_3(TPU_io_out_result_1_3),
    .io_out_cal(TPU_io_out_cal)
  );
  TPU TPU_1 ( // @[STA_VDBB.scala 97:36:@8677.4]
    .clock(TPU_1_clock),
    .reset(TPU_1_reset),
    .io_in_A_0_0(TPU_1_io_in_A_0_0),
    .io_in_A_0_1(TPU_1_io_in_A_0_1),
    .io_in_A_0_2(TPU_1_io_in_A_0_2),
    .io_in_A_0_3(TPU_1_io_in_A_0_3),
    .io_in_A_0_4(TPU_1_io_in_A_0_4),
    .io_in_A_0_5(TPU_1_io_in_A_0_5),
    .io_in_A_0_6(TPU_1_io_in_A_0_6),
    .io_in_A_0_7(TPU_1_io_in_A_0_7),
    .io_in_A_1_0(TPU_1_io_in_A_1_0),
    .io_in_A_1_1(TPU_1_io_in_A_1_1),
    .io_in_A_1_2(TPU_1_io_in_A_1_2),
    .io_in_A_1_3(TPU_1_io_in_A_1_3),
    .io_in_A_1_4(TPU_1_io_in_A_1_4),
    .io_in_A_1_5(TPU_1_io_in_A_1_5),
    .io_in_A_1_6(TPU_1_io_in_A_1_6),
    .io_in_A_1_7(TPU_1_io_in_A_1_7),
    .io_in_B_0_0(TPU_1_io_in_B_0_0),
    .io_in_B_0_1(TPU_1_io_in_B_0_1),
    .io_in_B_0_2(TPU_1_io_in_B_0_2),
    .io_in_B_0_3(TPU_1_io_in_B_0_3),
    .io_in_B_0_4(TPU_1_io_in_B_0_4),
    .io_in_B_0_5(TPU_1_io_in_B_0_5),
    .io_in_B_0_6(TPU_1_io_in_B_0_6),
    .io_in_B_0_7(TPU_1_io_in_B_0_7),
    .io_in_B_1_0(TPU_1_io_in_B_1_0),
    .io_in_B_1_1(TPU_1_io_in_B_1_1),
    .io_in_B_1_2(TPU_1_io_in_B_1_2),
    .io_in_B_1_3(TPU_1_io_in_B_1_3),
    .io_in_B_1_4(TPU_1_io_in_B_1_4),
    .io_in_B_1_5(TPU_1_io_in_B_1_5),
    .io_in_B_1_6(TPU_1_io_in_B_1_6),
    .io_in_B_1_7(TPU_1_io_in_B_1_7),
    .io_in_B_2_0(TPU_1_io_in_B_2_0),
    .io_in_B_2_1(TPU_1_io_in_B_2_1),
    .io_in_B_2_2(TPU_1_io_in_B_2_2),
    .io_in_B_2_3(TPU_1_io_in_B_2_3),
    .io_in_B_2_4(TPU_1_io_in_B_2_4),
    .io_in_B_2_5(TPU_1_io_in_B_2_5),
    .io_in_B_2_6(TPU_1_io_in_B_2_6),
    .io_in_B_2_7(TPU_1_io_in_B_2_7),
    .io_in_B_3_0(TPU_1_io_in_B_3_0),
    .io_in_B_3_1(TPU_1_io_in_B_3_1),
    .io_in_B_3_2(TPU_1_io_in_B_3_2),
    .io_in_B_3_3(TPU_1_io_in_B_3_3),
    .io_in_B_3_4(TPU_1_io_in_B_3_4),
    .io_in_B_3_5(TPU_1_io_in_B_3_5),
    .io_in_B_3_6(TPU_1_io_in_B_3_6),
    .io_in_B_3_7(TPU_1_io_in_B_3_7),
    .io_in_tag_0_0(TPU_1_io_in_tag_0_0),
    .io_in_tag_0_1(TPU_1_io_in_tag_0_1),
    .io_in_tag_0_2(TPU_1_io_in_tag_0_2),
    .io_in_tag_0_3(TPU_1_io_in_tag_0_3),
    .io_in_tag_0_4(TPU_1_io_in_tag_0_4),
    .io_in_tag_0_5(TPU_1_io_in_tag_0_5),
    .io_in_tag_0_6(TPU_1_io_in_tag_0_6),
    .io_in_tag_0_7(TPU_1_io_in_tag_0_7),
    .io_in_tag_1_0(TPU_1_io_in_tag_1_0),
    .io_in_tag_1_1(TPU_1_io_in_tag_1_1),
    .io_in_tag_1_2(TPU_1_io_in_tag_1_2),
    .io_in_tag_1_3(TPU_1_io_in_tag_1_3),
    .io_in_tag_1_4(TPU_1_io_in_tag_1_4),
    .io_in_tag_1_5(TPU_1_io_in_tag_1_5),
    .io_in_tag_1_6(TPU_1_io_in_tag_1_6),
    .io_in_tag_1_7(TPU_1_io_in_tag_1_7),
    .io_in_tag_2_0(TPU_1_io_in_tag_2_0),
    .io_in_tag_2_1(TPU_1_io_in_tag_2_1),
    .io_in_tag_2_2(TPU_1_io_in_tag_2_2),
    .io_in_tag_2_3(TPU_1_io_in_tag_2_3),
    .io_in_tag_2_4(TPU_1_io_in_tag_2_4),
    .io_in_tag_2_5(TPU_1_io_in_tag_2_5),
    .io_in_tag_2_6(TPU_1_io_in_tag_2_6),
    .io_in_tag_2_7(TPU_1_io_in_tag_2_7),
    .io_in_tag_3_0(TPU_1_io_in_tag_3_0),
    .io_in_tag_3_1(TPU_1_io_in_tag_3_1),
    .io_in_tag_3_2(TPU_1_io_in_tag_3_2),
    .io_in_tag_3_3(TPU_1_io_in_tag_3_3),
    .io_in_tag_3_4(TPU_1_io_in_tag_3_4),
    .io_in_tag_3_5(TPU_1_io_in_tag_3_5),
    .io_in_tag_3_6(TPU_1_io_in_tag_3_6),
    .io_in_tag_3_7(TPU_1_io_in_tag_3_7),
    .io_in_cal(TPU_1_io_in_cal),
    .io_out_A_0_0(TPU_1_io_out_A_0_0),
    .io_out_A_0_1(TPU_1_io_out_A_0_1),
    .io_out_A_0_2(TPU_1_io_out_A_0_2),
    .io_out_A_0_3(TPU_1_io_out_A_0_3),
    .io_out_A_0_4(TPU_1_io_out_A_0_4),
    .io_out_A_0_5(TPU_1_io_out_A_0_5),
    .io_out_A_0_6(TPU_1_io_out_A_0_6),
    .io_out_A_0_7(TPU_1_io_out_A_0_7),
    .io_out_A_1_0(TPU_1_io_out_A_1_0),
    .io_out_A_1_1(TPU_1_io_out_A_1_1),
    .io_out_A_1_2(TPU_1_io_out_A_1_2),
    .io_out_A_1_3(TPU_1_io_out_A_1_3),
    .io_out_A_1_4(TPU_1_io_out_A_1_4),
    .io_out_A_1_5(TPU_1_io_out_A_1_5),
    .io_out_A_1_6(TPU_1_io_out_A_1_6),
    .io_out_A_1_7(TPU_1_io_out_A_1_7),
    .io_out_B_0_0(TPU_1_io_out_B_0_0),
    .io_out_B_0_1(TPU_1_io_out_B_0_1),
    .io_out_B_0_2(TPU_1_io_out_B_0_2),
    .io_out_B_0_3(TPU_1_io_out_B_0_3),
    .io_out_B_0_4(TPU_1_io_out_B_0_4),
    .io_out_B_0_5(TPU_1_io_out_B_0_5),
    .io_out_B_0_6(TPU_1_io_out_B_0_6),
    .io_out_B_0_7(TPU_1_io_out_B_0_7),
    .io_out_B_1_0(TPU_1_io_out_B_1_0),
    .io_out_B_1_1(TPU_1_io_out_B_1_1),
    .io_out_B_1_2(TPU_1_io_out_B_1_2),
    .io_out_B_1_3(TPU_1_io_out_B_1_3),
    .io_out_B_1_4(TPU_1_io_out_B_1_4),
    .io_out_B_1_5(TPU_1_io_out_B_1_5),
    .io_out_B_1_6(TPU_1_io_out_B_1_6),
    .io_out_B_1_7(TPU_1_io_out_B_1_7),
    .io_out_B_2_0(TPU_1_io_out_B_2_0),
    .io_out_B_2_1(TPU_1_io_out_B_2_1),
    .io_out_B_2_2(TPU_1_io_out_B_2_2),
    .io_out_B_2_3(TPU_1_io_out_B_2_3),
    .io_out_B_2_4(TPU_1_io_out_B_2_4),
    .io_out_B_2_5(TPU_1_io_out_B_2_5),
    .io_out_B_2_6(TPU_1_io_out_B_2_6),
    .io_out_B_2_7(TPU_1_io_out_B_2_7),
    .io_out_B_3_0(TPU_1_io_out_B_3_0),
    .io_out_B_3_1(TPU_1_io_out_B_3_1),
    .io_out_B_3_2(TPU_1_io_out_B_3_2),
    .io_out_B_3_3(TPU_1_io_out_B_3_3),
    .io_out_B_3_4(TPU_1_io_out_B_3_4),
    .io_out_B_3_5(TPU_1_io_out_B_3_5),
    .io_out_B_3_6(TPU_1_io_out_B_3_6),
    .io_out_B_3_7(TPU_1_io_out_B_3_7),
    .io_out_tag_0_0(TPU_1_io_out_tag_0_0),
    .io_out_tag_0_1(TPU_1_io_out_tag_0_1),
    .io_out_tag_0_2(TPU_1_io_out_tag_0_2),
    .io_out_tag_0_3(TPU_1_io_out_tag_0_3),
    .io_out_tag_0_4(TPU_1_io_out_tag_0_4),
    .io_out_tag_0_5(TPU_1_io_out_tag_0_5),
    .io_out_tag_0_6(TPU_1_io_out_tag_0_6),
    .io_out_tag_0_7(TPU_1_io_out_tag_0_7),
    .io_out_tag_1_0(TPU_1_io_out_tag_1_0),
    .io_out_tag_1_1(TPU_1_io_out_tag_1_1),
    .io_out_tag_1_2(TPU_1_io_out_tag_1_2),
    .io_out_tag_1_3(TPU_1_io_out_tag_1_3),
    .io_out_tag_1_4(TPU_1_io_out_tag_1_4),
    .io_out_tag_1_5(TPU_1_io_out_tag_1_5),
    .io_out_tag_1_6(TPU_1_io_out_tag_1_6),
    .io_out_tag_1_7(TPU_1_io_out_tag_1_7),
    .io_out_tag_2_0(TPU_1_io_out_tag_2_0),
    .io_out_tag_2_1(TPU_1_io_out_tag_2_1),
    .io_out_tag_2_2(TPU_1_io_out_tag_2_2),
    .io_out_tag_2_3(TPU_1_io_out_tag_2_3),
    .io_out_tag_2_4(TPU_1_io_out_tag_2_4),
    .io_out_tag_2_5(TPU_1_io_out_tag_2_5),
    .io_out_tag_2_6(TPU_1_io_out_tag_2_6),
    .io_out_tag_2_7(TPU_1_io_out_tag_2_7),
    .io_out_tag_3_0(TPU_1_io_out_tag_3_0),
    .io_out_tag_3_1(TPU_1_io_out_tag_3_1),
    .io_out_tag_3_2(TPU_1_io_out_tag_3_2),
    .io_out_tag_3_3(TPU_1_io_out_tag_3_3),
    .io_out_tag_3_4(TPU_1_io_out_tag_3_4),
    .io_out_tag_3_5(TPU_1_io_out_tag_3_5),
    .io_out_tag_3_6(TPU_1_io_out_tag_3_6),
    .io_out_tag_3_7(TPU_1_io_out_tag_3_7),
    .io_out_result_0_0(TPU_1_io_out_result_0_0),
    .io_out_result_0_1(TPU_1_io_out_result_0_1),
    .io_out_result_0_2(TPU_1_io_out_result_0_2),
    .io_out_result_0_3(TPU_1_io_out_result_0_3),
    .io_out_result_1_0(TPU_1_io_out_result_1_0),
    .io_out_result_1_1(TPU_1_io_out_result_1_1),
    .io_out_result_1_2(TPU_1_io_out_result_1_2),
    .io_out_result_1_3(TPU_1_io_out_result_1_3),
    .io_out_cal(TPU_1_io_out_cal)
  );
  TPU TPU_2 ( // @[STA_VDBB.scala 97:36:@8680.4]
    .clock(TPU_2_clock),
    .reset(TPU_2_reset),
    .io_in_A_0_0(TPU_2_io_in_A_0_0),
    .io_in_A_0_1(TPU_2_io_in_A_0_1),
    .io_in_A_0_2(TPU_2_io_in_A_0_2),
    .io_in_A_0_3(TPU_2_io_in_A_0_3),
    .io_in_A_0_4(TPU_2_io_in_A_0_4),
    .io_in_A_0_5(TPU_2_io_in_A_0_5),
    .io_in_A_0_6(TPU_2_io_in_A_0_6),
    .io_in_A_0_7(TPU_2_io_in_A_0_7),
    .io_in_A_1_0(TPU_2_io_in_A_1_0),
    .io_in_A_1_1(TPU_2_io_in_A_1_1),
    .io_in_A_1_2(TPU_2_io_in_A_1_2),
    .io_in_A_1_3(TPU_2_io_in_A_1_3),
    .io_in_A_1_4(TPU_2_io_in_A_1_4),
    .io_in_A_1_5(TPU_2_io_in_A_1_5),
    .io_in_A_1_6(TPU_2_io_in_A_1_6),
    .io_in_A_1_7(TPU_2_io_in_A_1_7),
    .io_in_B_0_0(TPU_2_io_in_B_0_0),
    .io_in_B_0_1(TPU_2_io_in_B_0_1),
    .io_in_B_0_2(TPU_2_io_in_B_0_2),
    .io_in_B_0_3(TPU_2_io_in_B_0_3),
    .io_in_B_0_4(TPU_2_io_in_B_0_4),
    .io_in_B_0_5(TPU_2_io_in_B_0_5),
    .io_in_B_0_6(TPU_2_io_in_B_0_6),
    .io_in_B_0_7(TPU_2_io_in_B_0_7),
    .io_in_B_1_0(TPU_2_io_in_B_1_0),
    .io_in_B_1_1(TPU_2_io_in_B_1_1),
    .io_in_B_1_2(TPU_2_io_in_B_1_2),
    .io_in_B_1_3(TPU_2_io_in_B_1_3),
    .io_in_B_1_4(TPU_2_io_in_B_1_4),
    .io_in_B_1_5(TPU_2_io_in_B_1_5),
    .io_in_B_1_6(TPU_2_io_in_B_1_6),
    .io_in_B_1_7(TPU_2_io_in_B_1_7),
    .io_in_B_2_0(TPU_2_io_in_B_2_0),
    .io_in_B_2_1(TPU_2_io_in_B_2_1),
    .io_in_B_2_2(TPU_2_io_in_B_2_2),
    .io_in_B_2_3(TPU_2_io_in_B_2_3),
    .io_in_B_2_4(TPU_2_io_in_B_2_4),
    .io_in_B_2_5(TPU_2_io_in_B_2_5),
    .io_in_B_2_6(TPU_2_io_in_B_2_6),
    .io_in_B_2_7(TPU_2_io_in_B_2_7),
    .io_in_B_3_0(TPU_2_io_in_B_3_0),
    .io_in_B_3_1(TPU_2_io_in_B_3_1),
    .io_in_B_3_2(TPU_2_io_in_B_3_2),
    .io_in_B_3_3(TPU_2_io_in_B_3_3),
    .io_in_B_3_4(TPU_2_io_in_B_3_4),
    .io_in_B_3_5(TPU_2_io_in_B_3_5),
    .io_in_B_3_6(TPU_2_io_in_B_3_6),
    .io_in_B_3_7(TPU_2_io_in_B_3_7),
    .io_in_tag_0_0(TPU_2_io_in_tag_0_0),
    .io_in_tag_0_1(TPU_2_io_in_tag_0_1),
    .io_in_tag_0_2(TPU_2_io_in_tag_0_2),
    .io_in_tag_0_3(TPU_2_io_in_tag_0_3),
    .io_in_tag_0_4(TPU_2_io_in_tag_0_4),
    .io_in_tag_0_5(TPU_2_io_in_tag_0_5),
    .io_in_tag_0_6(TPU_2_io_in_tag_0_6),
    .io_in_tag_0_7(TPU_2_io_in_tag_0_7),
    .io_in_tag_1_0(TPU_2_io_in_tag_1_0),
    .io_in_tag_1_1(TPU_2_io_in_tag_1_1),
    .io_in_tag_1_2(TPU_2_io_in_tag_1_2),
    .io_in_tag_1_3(TPU_2_io_in_tag_1_3),
    .io_in_tag_1_4(TPU_2_io_in_tag_1_4),
    .io_in_tag_1_5(TPU_2_io_in_tag_1_5),
    .io_in_tag_1_6(TPU_2_io_in_tag_1_6),
    .io_in_tag_1_7(TPU_2_io_in_tag_1_7),
    .io_in_tag_2_0(TPU_2_io_in_tag_2_0),
    .io_in_tag_2_1(TPU_2_io_in_tag_2_1),
    .io_in_tag_2_2(TPU_2_io_in_tag_2_2),
    .io_in_tag_2_3(TPU_2_io_in_tag_2_3),
    .io_in_tag_2_4(TPU_2_io_in_tag_2_4),
    .io_in_tag_2_5(TPU_2_io_in_tag_2_5),
    .io_in_tag_2_6(TPU_2_io_in_tag_2_6),
    .io_in_tag_2_7(TPU_2_io_in_tag_2_7),
    .io_in_tag_3_0(TPU_2_io_in_tag_3_0),
    .io_in_tag_3_1(TPU_2_io_in_tag_3_1),
    .io_in_tag_3_2(TPU_2_io_in_tag_3_2),
    .io_in_tag_3_3(TPU_2_io_in_tag_3_3),
    .io_in_tag_3_4(TPU_2_io_in_tag_3_4),
    .io_in_tag_3_5(TPU_2_io_in_tag_3_5),
    .io_in_tag_3_6(TPU_2_io_in_tag_3_6),
    .io_in_tag_3_7(TPU_2_io_in_tag_3_7),
    .io_in_cal(TPU_2_io_in_cal),
    .io_out_A_0_0(TPU_2_io_out_A_0_0),
    .io_out_A_0_1(TPU_2_io_out_A_0_1),
    .io_out_A_0_2(TPU_2_io_out_A_0_2),
    .io_out_A_0_3(TPU_2_io_out_A_0_3),
    .io_out_A_0_4(TPU_2_io_out_A_0_4),
    .io_out_A_0_5(TPU_2_io_out_A_0_5),
    .io_out_A_0_6(TPU_2_io_out_A_0_6),
    .io_out_A_0_7(TPU_2_io_out_A_0_7),
    .io_out_A_1_0(TPU_2_io_out_A_1_0),
    .io_out_A_1_1(TPU_2_io_out_A_1_1),
    .io_out_A_1_2(TPU_2_io_out_A_1_2),
    .io_out_A_1_3(TPU_2_io_out_A_1_3),
    .io_out_A_1_4(TPU_2_io_out_A_1_4),
    .io_out_A_1_5(TPU_2_io_out_A_1_5),
    .io_out_A_1_6(TPU_2_io_out_A_1_6),
    .io_out_A_1_7(TPU_2_io_out_A_1_7),
    .io_out_B_0_0(TPU_2_io_out_B_0_0),
    .io_out_B_0_1(TPU_2_io_out_B_0_1),
    .io_out_B_0_2(TPU_2_io_out_B_0_2),
    .io_out_B_0_3(TPU_2_io_out_B_0_3),
    .io_out_B_0_4(TPU_2_io_out_B_0_4),
    .io_out_B_0_5(TPU_2_io_out_B_0_5),
    .io_out_B_0_6(TPU_2_io_out_B_0_6),
    .io_out_B_0_7(TPU_2_io_out_B_0_7),
    .io_out_B_1_0(TPU_2_io_out_B_1_0),
    .io_out_B_1_1(TPU_2_io_out_B_1_1),
    .io_out_B_1_2(TPU_2_io_out_B_1_2),
    .io_out_B_1_3(TPU_2_io_out_B_1_3),
    .io_out_B_1_4(TPU_2_io_out_B_1_4),
    .io_out_B_1_5(TPU_2_io_out_B_1_5),
    .io_out_B_1_6(TPU_2_io_out_B_1_6),
    .io_out_B_1_7(TPU_2_io_out_B_1_7),
    .io_out_B_2_0(TPU_2_io_out_B_2_0),
    .io_out_B_2_1(TPU_2_io_out_B_2_1),
    .io_out_B_2_2(TPU_2_io_out_B_2_2),
    .io_out_B_2_3(TPU_2_io_out_B_2_3),
    .io_out_B_2_4(TPU_2_io_out_B_2_4),
    .io_out_B_2_5(TPU_2_io_out_B_2_5),
    .io_out_B_2_6(TPU_2_io_out_B_2_6),
    .io_out_B_2_7(TPU_2_io_out_B_2_7),
    .io_out_B_3_0(TPU_2_io_out_B_3_0),
    .io_out_B_3_1(TPU_2_io_out_B_3_1),
    .io_out_B_3_2(TPU_2_io_out_B_3_2),
    .io_out_B_3_3(TPU_2_io_out_B_3_3),
    .io_out_B_3_4(TPU_2_io_out_B_3_4),
    .io_out_B_3_5(TPU_2_io_out_B_3_5),
    .io_out_B_3_6(TPU_2_io_out_B_3_6),
    .io_out_B_3_7(TPU_2_io_out_B_3_7),
    .io_out_tag_0_0(TPU_2_io_out_tag_0_0),
    .io_out_tag_0_1(TPU_2_io_out_tag_0_1),
    .io_out_tag_0_2(TPU_2_io_out_tag_0_2),
    .io_out_tag_0_3(TPU_2_io_out_tag_0_3),
    .io_out_tag_0_4(TPU_2_io_out_tag_0_4),
    .io_out_tag_0_5(TPU_2_io_out_tag_0_5),
    .io_out_tag_0_6(TPU_2_io_out_tag_0_6),
    .io_out_tag_0_7(TPU_2_io_out_tag_0_7),
    .io_out_tag_1_0(TPU_2_io_out_tag_1_0),
    .io_out_tag_1_1(TPU_2_io_out_tag_1_1),
    .io_out_tag_1_2(TPU_2_io_out_tag_1_2),
    .io_out_tag_1_3(TPU_2_io_out_tag_1_3),
    .io_out_tag_1_4(TPU_2_io_out_tag_1_4),
    .io_out_tag_1_5(TPU_2_io_out_tag_1_5),
    .io_out_tag_1_6(TPU_2_io_out_tag_1_6),
    .io_out_tag_1_7(TPU_2_io_out_tag_1_7),
    .io_out_tag_2_0(TPU_2_io_out_tag_2_0),
    .io_out_tag_2_1(TPU_2_io_out_tag_2_1),
    .io_out_tag_2_2(TPU_2_io_out_tag_2_2),
    .io_out_tag_2_3(TPU_2_io_out_tag_2_3),
    .io_out_tag_2_4(TPU_2_io_out_tag_2_4),
    .io_out_tag_2_5(TPU_2_io_out_tag_2_5),
    .io_out_tag_2_6(TPU_2_io_out_tag_2_6),
    .io_out_tag_2_7(TPU_2_io_out_tag_2_7),
    .io_out_tag_3_0(TPU_2_io_out_tag_3_0),
    .io_out_tag_3_1(TPU_2_io_out_tag_3_1),
    .io_out_tag_3_2(TPU_2_io_out_tag_3_2),
    .io_out_tag_3_3(TPU_2_io_out_tag_3_3),
    .io_out_tag_3_4(TPU_2_io_out_tag_3_4),
    .io_out_tag_3_5(TPU_2_io_out_tag_3_5),
    .io_out_tag_3_6(TPU_2_io_out_tag_3_6),
    .io_out_tag_3_7(TPU_2_io_out_tag_3_7),
    .io_out_result_0_0(TPU_2_io_out_result_0_0),
    .io_out_result_0_1(TPU_2_io_out_result_0_1),
    .io_out_result_0_2(TPU_2_io_out_result_0_2),
    .io_out_result_0_3(TPU_2_io_out_result_0_3),
    .io_out_result_1_0(TPU_2_io_out_result_1_0),
    .io_out_result_1_1(TPU_2_io_out_result_1_1),
    .io_out_result_1_2(TPU_2_io_out_result_1_2),
    .io_out_result_1_3(TPU_2_io_out_result_1_3),
    .io_out_cal(TPU_2_io_out_cal)
  );
  TPU TPU_3 ( // @[STA_VDBB.scala 97:36:@8683.4]
    .clock(TPU_3_clock),
    .reset(TPU_3_reset),
    .io_in_A_0_0(TPU_3_io_in_A_0_0),
    .io_in_A_0_1(TPU_3_io_in_A_0_1),
    .io_in_A_0_2(TPU_3_io_in_A_0_2),
    .io_in_A_0_3(TPU_3_io_in_A_0_3),
    .io_in_A_0_4(TPU_3_io_in_A_0_4),
    .io_in_A_0_5(TPU_3_io_in_A_0_5),
    .io_in_A_0_6(TPU_3_io_in_A_0_6),
    .io_in_A_0_7(TPU_3_io_in_A_0_7),
    .io_in_A_1_0(TPU_3_io_in_A_1_0),
    .io_in_A_1_1(TPU_3_io_in_A_1_1),
    .io_in_A_1_2(TPU_3_io_in_A_1_2),
    .io_in_A_1_3(TPU_3_io_in_A_1_3),
    .io_in_A_1_4(TPU_3_io_in_A_1_4),
    .io_in_A_1_5(TPU_3_io_in_A_1_5),
    .io_in_A_1_6(TPU_3_io_in_A_1_6),
    .io_in_A_1_7(TPU_3_io_in_A_1_7),
    .io_in_B_0_0(TPU_3_io_in_B_0_0),
    .io_in_B_0_1(TPU_3_io_in_B_0_1),
    .io_in_B_0_2(TPU_3_io_in_B_0_2),
    .io_in_B_0_3(TPU_3_io_in_B_0_3),
    .io_in_B_0_4(TPU_3_io_in_B_0_4),
    .io_in_B_0_5(TPU_3_io_in_B_0_5),
    .io_in_B_0_6(TPU_3_io_in_B_0_6),
    .io_in_B_0_7(TPU_3_io_in_B_0_7),
    .io_in_B_1_0(TPU_3_io_in_B_1_0),
    .io_in_B_1_1(TPU_3_io_in_B_1_1),
    .io_in_B_1_2(TPU_3_io_in_B_1_2),
    .io_in_B_1_3(TPU_3_io_in_B_1_3),
    .io_in_B_1_4(TPU_3_io_in_B_1_4),
    .io_in_B_1_5(TPU_3_io_in_B_1_5),
    .io_in_B_1_6(TPU_3_io_in_B_1_6),
    .io_in_B_1_7(TPU_3_io_in_B_1_7),
    .io_in_B_2_0(TPU_3_io_in_B_2_0),
    .io_in_B_2_1(TPU_3_io_in_B_2_1),
    .io_in_B_2_2(TPU_3_io_in_B_2_2),
    .io_in_B_2_3(TPU_3_io_in_B_2_3),
    .io_in_B_2_4(TPU_3_io_in_B_2_4),
    .io_in_B_2_5(TPU_3_io_in_B_2_5),
    .io_in_B_2_6(TPU_3_io_in_B_2_6),
    .io_in_B_2_7(TPU_3_io_in_B_2_7),
    .io_in_B_3_0(TPU_3_io_in_B_3_0),
    .io_in_B_3_1(TPU_3_io_in_B_3_1),
    .io_in_B_3_2(TPU_3_io_in_B_3_2),
    .io_in_B_3_3(TPU_3_io_in_B_3_3),
    .io_in_B_3_4(TPU_3_io_in_B_3_4),
    .io_in_B_3_5(TPU_3_io_in_B_3_5),
    .io_in_B_3_6(TPU_3_io_in_B_3_6),
    .io_in_B_3_7(TPU_3_io_in_B_3_7),
    .io_in_tag_0_0(TPU_3_io_in_tag_0_0),
    .io_in_tag_0_1(TPU_3_io_in_tag_0_1),
    .io_in_tag_0_2(TPU_3_io_in_tag_0_2),
    .io_in_tag_0_3(TPU_3_io_in_tag_0_3),
    .io_in_tag_0_4(TPU_3_io_in_tag_0_4),
    .io_in_tag_0_5(TPU_3_io_in_tag_0_5),
    .io_in_tag_0_6(TPU_3_io_in_tag_0_6),
    .io_in_tag_0_7(TPU_3_io_in_tag_0_7),
    .io_in_tag_1_0(TPU_3_io_in_tag_1_0),
    .io_in_tag_1_1(TPU_3_io_in_tag_1_1),
    .io_in_tag_1_2(TPU_3_io_in_tag_1_2),
    .io_in_tag_1_3(TPU_3_io_in_tag_1_3),
    .io_in_tag_1_4(TPU_3_io_in_tag_1_4),
    .io_in_tag_1_5(TPU_3_io_in_tag_1_5),
    .io_in_tag_1_6(TPU_3_io_in_tag_1_6),
    .io_in_tag_1_7(TPU_3_io_in_tag_1_7),
    .io_in_tag_2_0(TPU_3_io_in_tag_2_0),
    .io_in_tag_2_1(TPU_3_io_in_tag_2_1),
    .io_in_tag_2_2(TPU_3_io_in_tag_2_2),
    .io_in_tag_2_3(TPU_3_io_in_tag_2_3),
    .io_in_tag_2_4(TPU_3_io_in_tag_2_4),
    .io_in_tag_2_5(TPU_3_io_in_tag_2_5),
    .io_in_tag_2_6(TPU_3_io_in_tag_2_6),
    .io_in_tag_2_7(TPU_3_io_in_tag_2_7),
    .io_in_tag_3_0(TPU_3_io_in_tag_3_0),
    .io_in_tag_3_1(TPU_3_io_in_tag_3_1),
    .io_in_tag_3_2(TPU_3_io_in_tag_3_2),
    .io_in_tag_3_3(TPU_3_io_in_tag_3_3),
    .io_in_tag_3_4(TPU_3_io_in_tag_3_4),
    .io_in_tag_3_5(TPU_3_io_in_tag_3_5),
    .io_in_tag_3_6(TPU_3_io_in_tag_3_6),
    .io_in_tag_3_7(TPU_3_io_in_tag_3_7),
    .io_in_cal(TPU_3_io_in_cal),
    .io_out_A_0_0(TPU_3_io_out_A_0_0),
    .io_out_A_0_1(TPU_3_io_out_A_0_1),
    .io_out_A_0_2(TPU_3_io_out_A_0_2),
    .io_out_A_0_3(TPU_3_io_out_A_0_3),
    .io_out_A_0_4(TPU_3_io_out_A_0_4),
    .io_out_A_0_5(TPU_3_io_out_A_0_5),
    .io_out_A_0_6(TPU_3_io_out_A_0_6),
    .io_out_A_0_7(TPU_3_io_out_A_0_7),
    .io_out_A_1_0(TPU_3_io_out_A_1_0),
    .io_out_A_1_1(TPU_3_io_out_A_1_1),
    .io_out_A_1_2(TPU_3_io_out_A_1_2),
    .io_out_A_1_3(TPU_3_io_out_A_1_3),
    .io_out_A_1_4(TPU_3_io_out_A_1_4),
    .io_out_A_1_5(TPU_3_io_out_A_1_5),
    .io_out_A_1_6(TPU_3_io_out_A_1_6),
    .io_out_A_1_7(TPU_3_io_out_A_1_7),
    .io_out_B_0_0(TPU_3_io_out_B_0_0),
    .io_out_B_0_1(TPU_3_io_out_B_0_1),
    .io_out_B_0_2(TPU_3_io_out_B_0_2),
    .io_out_B_0_3(TPU_3_io_out_B_0_3),
    .io_out_B_0_4(TPU_3_io_out_B_0_4),
    .io_out_B_0_5(TPU_3_io_out_B_0_5),
    .io_out_B_0_6(TPU_3_io_out_B_0_6),
    .io_out_B_0_7(TPU_3_io_out_B_0_7),
    .io_out_B_1_0(TPU_3_io_out_B_1_0),
    .io_out_B_1_1(TPU_3_io_out_B_1_1),
    .io_out_B_1_2(TPU_3_io_out_B_1_2),
    .io_out_B_1_3(TPU_3_io_out_B_1_3),
    .io_out_B_1_4(TPU_3_io_out_B_1_4),
    .io_out_B_1_5(TPU_3_io_out_B_1_5),
    .io_out_B_1_6(TPU_3_io_out_B_1_6),
    .io_out_B_1_7(TPU_3_io_out_B_1_7),
    .io_out_B_2_0(TPU_3_io_out_B_2_0),
    .io_out_B_2_1(TPU_3_io_out_B_2_1),
    .io_out_B_2_2(TPU_3_io_out_B_2_2),
    .io_out_B_2_3(TPU_3_io_out_B_2_3),
    .io_out_B_2_4(TPU_3_io_out_B_2_4),
    .io_out_B_2_5(TPU_3_io_out_B_2_5),
    .io_out_B_2_6(TPU_3_io_out_B_2_6),
    .io_out_B_2_7(TPU_3_io_out_B_2_7),
    .io_out_B_3_0(TPU_3_io_out_B_3_0),
    .io_out_B_3_1(TPU_3_io_out_B_3_1),
    .io_out_B_3_2(TPU_3_io_out_B_3_2),
    .io_out_B_3_3(TPU_3_io_out_B_3_3),
    .io_out_B_3_4(TPU_3_io_out_B_3_4),
    .io_out_B_3_5(TPU_3_io_out_B_3_5),
    .io_out_B_3_6(TPU_3_io_out_B_3_6),
    .io_out_B_3_7(TPU_3_io_out_B_3_7),
    .io_out_tag_0_0(TPU_3_io_out_tag_0_0),
    .io_out_tag_0_1(TPU_3_io_out_tag_0_1),
    .io_out_tag_0_2(TPU_3_io_out_tag_0_2),
    .io_out_tag_0_3(TPU_3_io_out_tag_0_3),
    .io_out_tag_0_4(TPU_3_io_out_tag_0_4),
    .io_out_tag_0_5(TPU_3_io_out_tag_0_5),
    .io_out_tag_0_6(TPU_3_io_out_tag_0_6),
    .io_out_tag_0_7(TPU_3_io_out_tag_0_7),
    .io_out_tag_1_0(TPU_3_io_out_tag_1_0),
    .io_out_tag_1_1(TPU_3_io_out_tag_1_1),
    .io_out_tag_1_2(TPU_3_io_out_tag_1_2),
    .io_out_tag_1_3(TPU_3_io_out_tag_1_3),
    .io_out_tag_1_4(TPU_3_io_out_tag_1_4),
    .io_out_tag_1_5(TPU_3_io_out_tag_1_5),
    .io_out_tag_1_6(TPU_3_io_out_tag_1_6),
    .io_out_tag_1_7(TPU_3_io_out_tag_1_7),
    .io_out_tag_2_0(TPU_3_io_out_tag_2_0),
    .io_out_tag_2_1(TPU_3_io_out_tag_2_1),
    .io_out_tag_2_2(TPU_3_io_out_tag_2_2),
    .io_out_tag_2_3(TPU_3_io_out_tag_2_3),
    .io_out_tag_2_4(TPU_3_io_out_tag_2_4),
    .io_out_tag_2_5(TPU_3_io_out_tag_2_5),
    .io_out_tag_2_6(TPU_3_io_out_tag_2_6),
    .io_out_tag_2_7(TPU_3_io_out_tag_2_7),
    .io_out_tag_3_0(TPU_3_io_out_tag_3_0),
    .io_out_tag_3_1(TPU_3_io_out_tag_3_1),
    .io_out_tag_3_2(TPU_3_io_out_tag_3_2),
    .io_out_tag_3_3(TPU_3_io_out_tag_3_3),
    .io_out_tag_3_4(TPU_3_io_out_tag_3_4),
    .io_out_tag_3_5(TPU_3_io_out_tag_3_5),
    .io_out_tag_3_6(TPU_3_io_out_tag_3_6),
    .io_out_tag_3_7(TPU_3_io_out_tag_3_7),
    .io_out_result_0_0(TPU_3_io_out_result_0_0),
    .io_out_result_0_1(TPU_3_io_out_result_0_1),
    .io_out_result_0_2(TPU_3_io_out_result_0_2),
    .io_out_result_0_3(TPU_3_io_out_result_0_3),
    .io_out_result_1_0(TPU_3_io_out_result_1_0),
    .io_out_result_1_1(TPU_3_io_out_result_1_1),
    .io_out_result_1_2(TPU_3_io_out_result_1_2),
    .io_out_result_1_3(TPU_3_io_out_result_1_3),
    .io_out_cal(TPU_3_io_out_cal)
  );
  assign TPUs_1_out_cal = TPU_1_io_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8857.4]
  assign TPUs_2_out_cal = TPU_2_io_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9027.4]
  assign _T_40965 = TPUs_1_out_cal & TPUs_2_out_cal; // @[STA_VDBB.scala 115:35:@9857.4]
  assign _T_40966 = cal_state_0 & cal_state_1; // @[STA_VDBB.scala 117:30:@9860.4]
  assign _T_43000 = 3'h0 == stateReg; // @[Conditional.scala 37:30:@10008.4]
  assign _T_43004 = _T_43002 == 1'h0; // @[STA_VDBB.scala 143:24:@10012.6]
  assign _T_43005 = io_in_cal & _T_43004; // @[STA_VDBB.scala 143:22:@10013.6]
  assign _GEN_0 = _T_43005 ? 3'h1 : stateReg; // @[STA_VDBB.scala 143:44:@10014.6]
  assign _T_43006 = 3'h1 == stateReg; // @[Conditional.scala 37:30:@10019.6]
  assign _T_43007 = 1'h0 == loop_reg; // @[Conditional.scala 37:30:@10021.8]
  assign _GEN_1 = cal_state_0 ? 1'h0 : 1'h1; // @[STA_VDBB.scala 159:29:@10141.12]
  assign _GEN_2 = cal_state_0 ? 3'h2 : stateReg; // @[STA_VDBB.scala 159:29:@10141.12]
  assign _GEN_3 = cal_state_0 ? 1'h0 : loop_reg; // @[STA_VDBB.scala 159:29:@10141.12]
  assign _GEN_4 = loop_reg ? _GEN_1 : cal_control_0; // @[Conditional.scala 39:67:@10139.10]
  assign _GEN_5 = loop_reg ? _GEN_2 : stateReg; // @[Conditional.scala 39:67:@10139.10]
  assign _GEN_6 = loop_reg ? _GEN_3 : loop_reg; // @[Conditional.scala 39:67:@10139.10]
  assign _GEN_7 = _T_43007 ? $signed(reg_A_1_0_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_8 = _T_43007 ? $signed(reg_A_1_0_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_9 = _T_43007 ? $signed(reg_A_1_0_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_10 = _T_43007 ? $signed(reg_A_1_0_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_11 = _T_43007 ? $signed(reg_A_1_0_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_12 = _T_43007 ? $signed(reg_A_1_0_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_13 = _T_43007 ? $signed(reg_A_1_0_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_14 = _T_43007 ? $signed(reg_A_1_0_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_15 = _T_43007 ? $signed(reg_A_1_1_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_16 = _T_43007 ? $signed(reg_A_1_1_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_17 = _T_43007 ? $signed(reg_A_1_1_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_18 = _T_43007 ? $signed(reg_A_1_1_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_19 = _T_43007 ? $signed(reg_A_1_1_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_20 = _T_43007 ? $signed(reg_A_1_1_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_21 = _T_43007 ? $signed(reg_A_1_1_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_22 = _T_43007 ? $signed(reg_A_1_1_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_23 = _T_43007 ? $signed(reg_B_1_0_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_24 = _T_43007 ? $signed(reg_B_1_0_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_25 = _T_43007 ? $signed(reg_B_1_0_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_26 = _T_43007 ? $signed(reg_B_1_0_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_27 = _T_43007 ? $signed(reg_B_1_0_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_28 = _T_43007 ? $signed(reg_B_1_0_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_29 = _T_43007 ? $signed(reg_B_1_0_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_30 = _T_43007 ? $signed(reg_B_1_0_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_31 = _T_43007 ? $signed(reg_B_1_1_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_32 = _T_43007 ? $signed(reg_B_1_1_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_33 = _T_43007 ? $signed(reg_B_1_1_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_34 = _T_43007 ? $signed(reg_B_1_1_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_35 = _T_43007 ? $signed(reg_B_1_1_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_36 = _T_43007 ? $signed(reg_B_1_1_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_37 = _T_43007 ? $signed(reg_B_1_1_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_38 = _T_43007 ? $signed(reg_B_1_1_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_39 = _T_43007 ? $signed(reg_B_1_2_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_40 = _T_43007 ? $signed(reg_B_1_2_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_41 = _T_43007 ? $signed(reg_B_1_2_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_42 = _T_43007 ? $signed(reg_B_1_2_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_43 = _T_43007 ? $signed(reg_B_1_2_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_44 = _T_43007 ? $signed(reg_B_1_2_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_45 = _T_43007 ? $signed(reg_B_1_2_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_46 = _T_43007 ? $signed(reg_B_1_2_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_47 = _T_43007 ? $signed(reg_B_1_3_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_48 = _T_43007 ? $signed(reg_B_1_3_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_49 = _T_43007 ? $signed(reg_B_1_3_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_50 = _T_43007 ? $signed(reg_B_1_3_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_51 = _T_43007 ? $signed(reg_B_1_3_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_52 = _T_43007 ? $signed(reg_B_1_3_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_53 = _T_43007 ? $signed(reg_B_1_3_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_54 = _T_43007 ? $signed(reg_B_1_3_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_119 = _T_43007 ? 1'h1 : _GEN_6; // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_120 = _T_43007 ? cal_control_0 : _GEN_4; // @[Conditional.scala 40:58:@10022.8]
  assign _GEN_121 = _T_43007 ? stateReg : _GEN_5; // @[Conditional.scala 40:58:@10022.8]
  assign _T_43011 = 3'h2 == stateReg; // @[Conditional.scala 37:30:@10149.8]
  assign _GEN_122 = cal_state_1 ? 1'h0 : 1'h1; // @[STA_VDBB.scala 179:29:@10271.14]
  assign _GEN_123 = cal_state_1 ? 3'h3 : stateReg; // @[STA_VDBB.scala 179:29:@10271.14]
  assign _GEN_124 = cal_state_1 ? 1'h0 : loop_reg; // @[STA_VDBB.scala 179:29:@10271.14]
  assign _GEN_125 = loop_reg ? _GEN_122 : cal_control_1; // @[Conditional.scala 39:67:@10269.12]
  assign _GEN_126 = loop_reg ? _GEN_123 : stateReg; // @[Conditional.scala 39:67:@10269.12]
  assign _GEN_127 = loop_reg ? _GEN_124 : loop_reg; // @[Conditional.scala 39:67:@10269.12]
  assign TPUs_0_out_A_0_0 = TPU_io_out_A_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8760.4]
  assign _GEN_128 = _T_43007 ? $signed(reg_A_2_0_0) : $signed(TPUs_0_out_A_0_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_1 = TPU_io_out_A_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8761.4]
  assign _GEN_129 = _T_43007 ? $signed(reg_A_2_0_1) : $signed(TPUs_0_out_A_0_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_2 = TPU_io_out_A_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8762.4]
  assign _GEN_130 = _T_43007 ? $signed(reg_A_2_0_2) : $signed(TPUs_0_out_A_0_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_3 = TPU_io_out_A_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8763.4]
  assign _GEN_131 = _T_43007 ? $signed(reg_A_2_0_3) : $signed(TPUs_0_out_A_0_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_4 = TPU_io_out_A_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8764.4]
  assign _GEN_132 = _T_43007 ? $signed(reg_A_2_0_4) : $signed(TPUs_0_out_A_0_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_5 = TPU_io_out_A_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8765.4]
  assign _GEN_133 = _T_43007 ? $signed(reg_A_2_0_5) : $signed(TPUs_0_out_A_0_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_6 = TPU_io_out_A_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8766.4]
  assign _GEN_134 = _T_43007 ? $signed(reg_A_2_0_6) : $signed(TPUs_0_out_A_0_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_0_7 = TPU_io_out_A_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8767.4]
  assign _GEN_135 = _T_43007 ? $signed(reg_A_2_0_7) : $signed(TPUs_0_out_A_0_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_0 = TPU_io_out_A_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8768.4]
  assign _GEN_136 = _T_43007 ? $signed(reg_A_2_1_0) : $signed(TPUs_0_out_A_1_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_1 = TPU_io_out_A_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8769.4]
  assign _GEN_137 = _T_43007 ? $signed(reg_A_2_1_1) : $signed(TPUs_0_out_A_1_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_2 = TPU_io_out_A_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8770.4]
  assign _GEN_138 = _T_43007 ? $signed(reg_A_2_1_2) : $signed(TPUs_0_out_A_1_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_3 = TPU_io_out_A_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8771.4]
  assign _GEN_139 = _T_43007 ? $signed(reg_A_2_1_3) : $signed(TPUs_0_out_A_1_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_4 = TPU_io_out_A_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8772.4]
  assign _GEN_140 = _T_43007 ? $signed(reg_A_2_1_4) : $signed(TPUs_0_out_A_1_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_5 = TPU_io_out_A_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8773.4]
  assign _GEN_141 = _T_43007 ? $signed(reg_A_2_1_5) : $signed(TPUs_0_out_A_1_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_6 = TPU_io_out_A_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8774.4]
  assign _GEN_142 = _T_43007 ? $signed(reg_A_2_1_6) : $signed(TPUs_0_out_A_1_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_A_1_7 = TPU_io_out_A_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8775.4]
  assign _GEN_143 = _T_43007 ? $signed(reg_A_2_1_7) : $signed(TPUs_0_out_A_1_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_0 = TPU_io_out_B_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8728.4]
  assign _GEN_144 = _T_43007 ? $signed(reg_B_2_0_0) : $signed(TPUs_0_out_B_0_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_1 = TPU_io_out_B_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8729.4]
  assign _GEN_145 = _T_43007 ? $signed(reg_B_2_0_1) : $signed(TPUs_0_out_B_0_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_2 = TPU_io_out_B_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8730.4]
  assign _GEN_146 = _T_43007 ? $signed(reg_B_2_0_2) : $signed(TPUs_0_out_B_0_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_3 = TPU_io_out_B_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8731.4]
  assign _GEN_147 = _T_43007 ? $signed(reg_B_2_0_3) : $signed(TPUs_0_out_B_0_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_4 = TPU_io_out_B_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8732.4]
  assign _GEN_148 = _T_43007 ? $signed(reg_B_2_0_4) : $signed(TPUs_0_out_B_0_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_5 = TPU_io_out_B_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8733.4]
  assign _GEN_149 = _T_43007 ? $signed(reg_B_2_0_5) : $signed(TPUs_0_out_B_0_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_6 = TPU_io_out_B_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8734.4]
  assign _GEN_150 = _T_43007 ? $signed(reg_B_2_0_6) : $signed(TPUs_0_out_B_0_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_0_7 = TPU_io_out_B_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8735.4]
  assign _GEN_151 = _T_43007 ? $signed(reg_B_2_0_7) : $signed(TPUs_0_out_B_0_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_0 = TPU_io_out_B_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8736.4]
  assign _GEN_152 = _T_43007 ? $signed(reg_B_2_1_0) : $signed(TPUs_0_out_B_1_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_1 = TPU_io_out_B_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8737.4]
  assign _GEN_153 = _T_43007 ? $signed(reg_B_2_1_1) : $signed(TPUs_0_out_B_1_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_2 = TPU_io_out_B_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8738.4]
  assign _GEN_154 = _T_43007 ? $signed(reg_B_2_1_2) : $signed(TPUs_0_out_B_1_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_3 = TPU_io_out_B_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8739.4]
  assign _GEN_155 = _T_43007 ? $signed(reg_B_2_1_3) : $signed(TPUs_0_out_B_1_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_4 = TPU_io_out_B_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8740.4]
  assign _GEN_156 = _T_43007 ? $signed(reg_B_2_1_4) : $signed(TPUs_0_out_B_1_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_5 = TPU_io_out_B_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8741.4]
  assign _GEN_157 = _T_43007 ? $signed(reg_B_2_1_5) : $signed(TPUs_0_out_B_1_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_6 = TPU_io_out_B_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8742.4]
  assign _GEN_158 = _T_43007 ? $signed(reg_B_2_1_6) : $signed(TPUs_0_out_B_1_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_1_7 = TPU_io_out_B_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8743.4]
  assign _GEN_159 = _T_43007 ? $signed(reg_B_2_1_7) : $signed(TPUs_0_out_B_1_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_0 = TPU_io_out_B_2_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8744.4]
  assign _GEN_160 = _T_43007 ? $signed(reg_B_2_2_0) : $signed(TPUs_0_out_B_2_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_1 = TPU_io_out_B_2_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8745.4]
  assign _GEN_161 = _T_43007 ? $signed(reg_B_2_2_1) : $signed(TPUs_0_out_B_2_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_2 = TPU_io_out_B_2_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8746.4]
  assign _GEN_162 = _T_43007 ? $signed(reg_B_2_2_2) : $signed(TPUs_0_out_B_2_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_3 = TPU_io_out_B_2_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8747.4]
  assign _GEN_163 = _T_43007 ? $signed(reg_B_2_2_3) : $signed(TPUs_0_out_B_2_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_4 = TPU_io_out_B_2_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8748.4]
  assign _GEN_164 = _T_43007 ? $signed(reg_B_2_2_4) : $signed(TPUs_0_out_B_2_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_5 = TPU_io_out_B_2_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8749.4]
  assign _GEN_165 = _T_43007 ? $signed(reg_B_2_2_5) : $signed(TPUs_0_out_B_2_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_6 = TPU_io_out_B_2_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8750.4]
  assign _GEN_166 = _T_43007 ? $signed(reg_B_2_2_6) : $signed(TPUs_0_out_B_2_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_2_7 = TPU_io_out_B_2_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8751.4]
  assign _GEN_167 = _T_43007 ? $signed(reg_B_2_2_7) : $signed(TPUs_0_out_B_2_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_0 = TPU_io_out_B_3_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8752.4]
  assign _GEN_168 = _T_43007 ? $signed(reg_B_2_3_0) : $signed(TPUs_0_out_B_3_0); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_1 = TPU_io_out_B_3_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8753.4]
  assign _GEN_169 = _T_43007 ? $signed(reg_B_2_3_1) : $signed(TPUs_0_out_B_3_1); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_2 = TPU_io_out_B_3_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8754.4]
  assign _GEN_170 = _T_43007 ? $signed(reg_B_2_3_2) : $signed(TPUs_0_out_B_3_2); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_3 = TPU_io_out_B_3_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8755.4]
  assign _GEN_171 = _T_43007 ? $signed(reg_B_2_3_3) : $signed(TPUs_0_out_B_3_3); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_4 = TPU_io_out_B_3_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8756.4]
  assign _GEN_172 = _T_43007 ? $signed(reg_B_2_3_4) : $signed(TPUs_0_out_B_3_4); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_5 = TPU_io_out_B_3_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8757.4]
  assign _GEN_173 = _T_43007 ? $signed(reg_B_2_3_5) : $signed(TPUs_0_out_B_3_5); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_6 = TPU_io_out_B_3_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8758.4]
  assign _GEN_174 = _T_43007 ? $signed(reg_B_2_3_6) : $signed(TPUs_0_out_B_3_6); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_B_3_7 = TPU_io_out_B_3_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8759.4]
  assign _GEN_175 = _T_43007 ? $signed(reg_B_2_3_7) : $signed(TPUs_0_out_B_3_7); // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_0 = TPU_io_out_tag_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8696.4]
  assign _GEN_208 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_0; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_1 = TPU_io_out_tag_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8697.4]
  assign _GEN_209 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_1; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_2 = TPU_io_out_tag_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8698.4]
  assign _GEN_210 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_2; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_3 = TPU_io_out_tag_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8699.4]
  assign _GEN_211 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_3; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_4 = TPU_io_out_tag_0_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8700.4]
  assign _GEN_212 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_4; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_5 = TPU_io_out_tag_0_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8701.4]
  assign _GEN_213 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_5; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_6 = TPU_io_out_tag_0_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8702.4]
  assign _GEN_214 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_6; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_0_7 = TPU_io_out_tag_0_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8703.4]
  assign _GEN_215 = _T_43007 ? 1'h0 : TPUs_0_out_tag_0_7; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_0 = TPU_io_out_tag_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8704.4]
  assign _GEN_216 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_0; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_1 = TPU_io_out_tag_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8705.4]
  assign _GEN_217 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_1; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_2 = TPU_io_out_tag_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8706.4]
  assign _GEN_218 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_2; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_3 = TPU_io_out_tag_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8707.4]
  assign _GEN_219 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_3; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_4 = TPU_io_out_tag_1_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8708.4]
  assign _GEN_220 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_4; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_5 = TPU_io_out_tag_1_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8709.4]
  assign _GEN_221 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_5; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_6 = TPU_io_out_tag_1_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8710.4]
  assign _GEN_222 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_6; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_1_7 = TPU_io_out_tag_1_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8711.4]
  assign _GEN_223 = _T_43007 ? 1'h0 : TPUs_0_out_tag_1_7; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_0 = TPU_io_out_tag_2_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8712.4]
  assign _GEN_224 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_0; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_1 = TPU_io_out_tag_2_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8713.4]
  assign _GEN_225 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_1; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_2 = TPU_io_out_tag_2_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8714.4]
  assign _GEN_226 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_2; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_3 = TPU_io_out_tag_2_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8715.4]
  assign _GEN_227 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_3; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_4 = TPU_io_out_tag_2_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8716.4]
  assign _GEN_228 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_4; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_5 = TPU_io_out_tag_2_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8717.4]
  assign _GEN_229 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_5; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_6 = TPU_io_out_tag_2_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8718.4]
  assign _GEN_230 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_6; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_2_7 = TPU_io_out_tag_2_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8719.4]
  assign _GEN_231 = _T_43007 ? 1'h0 : TPUs_0_out_tag_2_7; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_0 = TPU_io_out_tag_3_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8720.4]
  assign _GEN_232 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_0; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_1 = TPU_io_out_tag_3_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8721.4]
  assign _GEN_233 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_1; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_2 = TPU_io_out_tag_3_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8722.4]
  assign _GEN_234 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_2; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_3 = TPU_io_out_tag_3_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8723.4]
  assign _GEN_235 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_3; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_4 = TPU_io_out_tag_3_4; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8724.4]
  assign _GEN_236 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_4; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_5 = TPU_io_out_tag_3_5; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8725.4]
  assign _GEN_237 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_5; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_6 = TPU_io_out_tag_3_6; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8726.4]
  assign _GEN_238 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_6; // @[Conditional.scala 40:58:@10152.10]
  assign TPUs_0_out_tag_3_7 = TPU_io_out_tag_3_7; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8727.4]
  assign _GEN_239 = _T_43007 ? 1'h0 : TPUs_0_out_tag_3_7; // @[Conditional.scala 40:58:@10152.10]
  assign _GEN_240 = _T_43007 ? 1'h1 : _GEN_127; // @[Conditional.scala 40:58:@10152.10]
  assign _GEN_241 = _T_43007 ? cal_control_1 : _GEN_125; // @[Conditional.scala 40:58:@10152.10]
  assign _GEN_242 = _T_43007 ? stateReg : _GEN_126; // @[Conditional.scala 40:58:@10152.10]
  assign _T_43016 = 3'h3 == stateReg; // @[Conditional.scala 37:30:@10279.10]
  assign _T_43021 = cal_state_0 & cal_state_2; // @[STA_VDBB.scala 200:29:@10402.16]
  assign _GEN_243 = _T_43021 ? 1'h0 : 1'h1; // @[STA_VDBB.scala 200:45:@10403.16]
  assign _GEN_244 = _T_43021 ? 3'h4 : stateReg; // @[STA_VDBB.scala 200:45:@10403.16]
  assign _GEN_245 = _T_43021 ? 1'h0 : loop_reg; // @[STA_VDBB.scala 200:45:@10403.16]
  assign _GEN_246 = loop_reg ? _GEN_243 : cal_control_0; // @[Conditional.scala 39:67:@10399.14]
  assign _GEN_247 = loop_reg ? _GEN_243 : cal_control_2; // @[Conditional.scala 39:67:@10399.14]
  assign _GEN_248 = loop_reg ? _GEN_244 : stateReg; // @[Conditional.scala 39:67:@10399.14]
  assign _GEN_249 = loop_reg ? _GEN_245 : loop_reg; // @[Conditional.scala 39:67:@10399.14]
  assign _GEN_250 = _T_43007 ? $signed(reg_A_3_0_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_251 = _T_43007 ? $signed(reg_A_3_0_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_252 = _T_43007 ? $signed(reg_A_3_0_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_253 = _T_43007 ? $signed(reg_A_3_0_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_254 = _T_43007 ? $signed(reg_A_3_0_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_255 = _T_43007 ? $signed(reg_A_3_0_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_256 = _T_43007 ? $signed(reg_A_3_0_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_257 = _T_43007 ? $signed(reg_A_3_0_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_258 = _T_43007 ? $signed(reg_A_3_1_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_259 = _T_43007 ? $signed(reg_A_3_1_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_260 = _T_43007 ? $signed(reg_A_3_1_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_261 = _T_43007 ? $signed(reg_A_3_1_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_262 = _T_43007 ? $signed(reg_A_3_1_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_263 = _T_43007 ? $signed(reg_A_3_1_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_264 = _T_43007 ? $signed(reg_A_3_1_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_265 = _T_43007 ? $signed(reg_A_3_1_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_266 = _T_43007 ? $signed(reg_B_3_0_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_267 = _T_43007 ? $signed(reg_B_3_0_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_268 = _T_43007 ? $signed(reg_B_3_0_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_269 = _T_43007 ? $signed(reg_B_3_0_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_270 = _T_43007 ? $signed(reg_B_3_0_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_271 = _T_43007 ? $signed(reg_B_3_0_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_272 = _T_43007 ? $signed(reg_B_3_0_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_273 = _T_43007 ? $signed(reg_B_3_0_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_274 = _T_43007 ? $signed(reg_B_3_1_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_275 = _T_43007 ? $signed(reg_B_3_1_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_276 = _T_43007 ? $signed(reg_B_3_1_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_277 = _T_43007 ? $signed(reg_B_3_1_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_278 = _T_43007 ? $signed(reg_B_3_1_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_279 = _T_43007 ? $signed(reg_B_3_1_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_280 = _T_43007 ? $signed(reg_B_3_1_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_281 = _T_43007 ? $signed(reg_B_3_1_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_282 = _T_43007 ? $signed(reg_B_3_2_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_283 = _T_43007 ? $signed(reg_B_3_2_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_284 = _T_43007 ? $signed(reg_B_3_2_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_285 = _T_43007 ? $signed(reg_B_3_2_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_286 = _T_43007 ? $signed(reg_B_3_2_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_287 = _T_43007 ? $signed(reg_B_3_2_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_288 = _T_43007 ? $signed(reg_B_3_2_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_289 = _T_43007 ? $signed(reg_B_3_2_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_290 = _T_43007 ? $signed(reg_B_3_3_0) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_291 = _T_43007 ? $signed(reg_B_3_3_1) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_292 = _T_43007 ? $signed(reg_B_3_3_2) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_293 = _T_43007 ? $signed(reg_B_3_3_3) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_294 = _T_43007 ? $signed(reg_B_3_3_4) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_295 = _T_43007 ? $signed(reg_B_3_3_5) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_296 = _T_43007 ? $signed(reg_B_3_3_6) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_297 = _T_43007 ? $signed(reg_B_3_3_7) : $signed(32'sh0); // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_362 = _T_43007 ? 1'h1 : _GEN_249; // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_363 = _T_43007 ? cal_control_0 : _GEN_246; // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_364 = _T_43007 ? cal_control_2 : _GEN_247; // @[Conditional.scala 40:58:@10282.12]
  assign _GEN_365 = _T_43007 ? stateReg : _GEN_248; // @[Conditional.scala 40:58:@10282.12]
  assign _T_43024 = 3'h4 == stateReg; // @[Conditional.scala 37:30:@10412.12]
  assign _GEN_366 = cal_state_1 ? 3'h5 : stateReg; // @[STA_VDBB.scala 221:29:@10534.18]
  assign _GEN_368 = loop_reg ? _GEN_366 : stateReg; // @[Conditional.scala 39:67:@10532.16]
  assign _GEN_370 = _T_43007 ? $signed(reg_A_4_0_0) : $signed(TPUs_0_out_A_0_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_371 = _T_43007 ? $signed(reg_A_4_0_1) : $signed(TPUs_0_out_A_0_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_372 = _T_43007 ? $signed(reg_A_4_0_2) : $signed(TPUs_0_out_A_0_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_373 = _T_43007 ? $signed(reg_A_4_0_3) : $signed(TPUs_0_out_A_0_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_374 = _T_43007 ? $signed(reg_A_4_0_4) : $signed(TPUs_0_out_A_0_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_375 = _T_43007 ? $signed(reg_A_4_0_5) : $signed(TPUs_0_out_A_0_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_376 = _T_43007 ? $signed(reg_A_4_0_6) : $signed(TPUs_0_out_A_0_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_377 = _T_43007 ? $signed(reg_A_4_0_7) : $signed(TPUs_0_out_A_0_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_378 = _T_43007 ? $signed(reg_A_4_1_0) : $signed(TPUs_0_out_A_1_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_379 = _T_43007 ? $signed(reg_A_4_1_1) : $signed(TPUs_0_out_A_1_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_380 = _T_43007 ? $signed(reg_A_4_1_2) : $signed(TPUs_0_out_A_1_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_381 = _T_43007 ? $signed(reg_A_4_1_3) : $signed(TPUs_0_out_A_1_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_382 = _T_43007 ? $signed(reg_A_4_1_4) : $signed(TPUs_0_out_A_1_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_383 = _T_43007 ? $signed(reg_A_4_1_5) : $signed(TPUs_0_out_A_1_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_384 = _T_43007 ? $signed(reg_A_4_1_6) : $signed(TPUs_0_out_A_1_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_385 = _T_43007 ? $signed(reg_A_4_1_7) : $signed(TPUs_0_out_A_1_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_386 = _T_43007 ? $signed(reg_B_4_0_0) : $signed(TPUs_0_out_B_0_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_387 = _T_43007 ? $signed(reg_B_4_0_1) : $signed(TPUs_0_out_B_0_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_388 = _T_43007 ? $signed(reg_B_4_0_2) : $signed(TPUs_0_out_B_0_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_389 = _T_43007 ? $signed(reg_B_4_0_3) : $signed(TPUs_0_out_B_0_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_390 = _T_43007 ? $signed(reg_B_4_0_4) : $signed(TPUs_0_out_B_0_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_391 = _T_43007 ? $signed(reg_B_4_0_5) : $signed(TPUs_0_out_B_0_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_392 = _T_43007 ? $signed(reg_B_4_0_6) : $signed(TPUs_0_out_B_0_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_393 = _T_43007 ? $signed(reg_B_4_0_7) : $signed(TPUs_0_out_B_0_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_394 = _T_43007 ? $signed(reg_B_4_1_0) : $signed(TPUs_0_out_B_1_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_395 = _T_43007 ? $signed(reg_B_4_1_1) : $signed(TPUs_0_out_B_1_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_396 = _T_43007 ? $signed(reg_B_4_1_2) : $signed(TPUs_0_out_B_1_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_397 = _T_43007 ? $signed(reg_B_4_1_3) : $signed(TPUs_0_out_B_1_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_398 = _T_43007 ? $signed(reg_B_4_1_4) : $signed(TPUs_0_out_B_1_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_399 = _T_43007 ? $signed(reg_B_4_1_5) : $signed(TPUs_0_out_B_1_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_400 = _T_43007 ? $signed(reg_B_4_1_6) : $signed(TPUs_0_out_B_1_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_401 = _T_43007 ? $signed(reg_B_4_1_7) : $signed(TPUs_0_out_B_1_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_402 = _T_43007 ? $signed(reg_B_4_2_0) : $signed(TPUs_0_out_B_2_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_403 = _T_43007 ? $signed(reg_B_4_2_1) : $signed(TPUs_0_out_B_2_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_404 = _T_43007 ? $signed(reg_B_4_2_2) : $signed(TPUs_0_out_B_2_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_405 = _T_43007 ? $signed(reg_B_4_2_3) : $signed(TPUs_0_out_B_2_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_406 = _T_43007 ? $signed(reg_B_4_2_4) : $signed(TPUs_0_out_B_2_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_407 = _T_43007 ? $signed(reg_B_4_2_5) : $signed(TPUs_0_out_B_2_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_408 = _T_43007 ? $signed(reg_B_4_2_6) : $signed(TPUs_0_out_B_2_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_409 = _T_43007 ? $signed(reg_B_4_2_7) : $signed(TPUs_0_out_B_2_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_410 = _T_43007 ? $signed(reg_B_4_3_0) : $signed(TPUs_0_out_B_3_0); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_411 = _T_43007 ? $signed(reg_B_4_3_1) : $signed(TPUs_0_out_B_3_1); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_412 = _T_43007 ? $signed(reg_B_4_3_2) : $signed(TPUs_0_out_B_3_2); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_413 = _T_43007 ? $signed(reg_B_4_3_3) : $signed(TPUs_0_out_B_3_3); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_414 = _T_43007 ? $signed(reg_B_4_3_4) : $signed(TPUs_0_out_B_3_4); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_415 = _T_43007 ? $signed(reg_B_4_3_5) : $signed(TPUs_0_out_B_3_5); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_416 = _T_43007 ? $signed(reg_B_4_3_6) : $signed(TPUs_0_out_B_3_6); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_417 = _T_43007 ? $signed(reg_B_4_3_7) : $signed(TPUs_0_out_B_3_7); // @[Conditional.scala 40:58:@10415.14]
  assign _GEN_484 = _T_43007 ? stateReg : _GEN_368; // @[Conditional.scala 40:58:@10415.14]
  assign _T_43029 = 3'h5 == stateReg; // @[Conditional.scala 37:30:@10542.14]
  assign _GEN_485 = cal_state_2 ? 1'h0 : cal_control_0; // @[STA_VDBB.scala 237:29:@10552.20]
  assign _GEN_486 = cal_state_2 ? 3'h0 : stateReg; // @[STA_VDBB.scala 237:29:@10552.20]
  assign _GEN_487 = cal_state_2 ? 1'h0 : loop_reg; // @[STA_VDBB.scala 237:29:@10552.20]
  assign _GEN_488 = loop_reg ? 1'h1 : cal_control_2; // @[Conditional.scala 39:67:@10550.18]
  assign _GEN_489 = loop_reg ? _GEN_485 : cal_control_0; // @[Conditional.scala 39:67:@10550.18]
  assign _GEN_490 = loop_reg ? _GEN_486 : stateReg; // @[Conditional.scala 39:67:@10550.18]
  assign _GEN_491 = loop_reg ? _GEN_487 : loop_reg; // @[Conditional.scala 39:67:@10550.18]
  assign _GEN_492 = _T_43007 ? 1'h1 : _GEN_491; // @[Conditional.scala 40:58:@10545.16]
  assign _GEN_493 = _T_43007 ? cal_control_2 : _GEN_488; // @[Conditional.scala 40:58:@10545.16]
  assign _GEN_494 = _T_43007 ? cal_control_0 : _GEN_489; // @[Conditional.scala 40:58:@10545.16]
  assign _GEN_495 = _T_43007 ? stateReg : _GEN_490; // @[Conditional.scala 40:58:@10545.16]
  assign _GEN_496 = _T_43029 ? _GEN_492 : loop_reg; // @[Conditional.scala 39:67:@10543.14]
  assign _GEN_497 = _T_43029 ? _GEN_493 : cal_control_2; // @[Conditional.scala 39:67:@10543.14]
  assign _GEN_498 = _T_43029 ? _GEN_494 : cal_control_0; // @[Conditional.scala 39:67:@10543.14]
  assign _GEN_499 = _T_43029 ? _GEN_495 : stateReg; // @[Conditional.scala 39:67:@10543.14]
  assign _GEN_500 = _T_43024 ? $signed(_GEN_370) : $signed(TPUs_0_out_A_0_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_501 = _T_43024 ? $signed(_GEN_371) : $signed(TPUs_0_out_A_0_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_502 = _T_43024 ? $signed(_GEN_372) : $signed(TPUs_0_out_A_0_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_503 = _T_43024 ? $signed(_GEN_373) : $signed(TPUs_0_out_A_0_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_504 = _T_43024 ? $signed(_GEN_374) : $signed(TPUs_0_out_A_0_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_505 = _T_43024 ? $signed(_GEN_375) : $signed(TPUs_0_out_A_0_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_506 = _T_43024 ? $signed(_GEN_376) : $signed(TPUs_0_out_A_0_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_507 = _T_43024 ? $signed(_GEN_377) : $signed(TPUs_0_out_A_0_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_508 = _T_43024 ? $signed(_GEN_378) : $signed(TPUs_0_out_A_1_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_509 = _T_43024 ? $signed(_GEN_379) : $signed(TPUs_0_out_A_1_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_510 = _T_43024 ? $signed(_GEN_380) : $signed(TPUs_0_out_A_1_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_511 = _T_43024 ? $signed(_GEN_381) : $signed(TPUs_0_out_A_1_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_512 = _T_43024 ? $signed(_GEN_382) : $signed(TPUs_0_out_A_1_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_513 = _T_43024 ? $signed(_GEN_383) : $signed(TPUs_0_out_A_1_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_514 = _T_43024 ? $signed(_GEN_384) : $signed(TPUs_0_out_A_1_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_515 = _T_43024 ? $signed(_GEN_385) : $signed(TPUs_0_out_A_1_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_516 = _T_43024 ? $signed(_GEN_386) : $signed(TPUs_0_out_B_0_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_517 = _T_43024 ? $signed(_GEN_387) : $signed(TPUs_0_out_B_0_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_518 = _T_43024 ? $signed(_GEN_388) : $signed(TPUs_0_out_B_0_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_519 = _T_43024 ? $signed(_GEN_389) : $signed(TPUs_0_out_B_0_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_520 = _T_43024 ? $signed(_GEN_390) : $signed(TPUs_0_out_B_0_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_521 = _T_43024 ? $signed(_GEN_391) : $signed(TPUs_0_out_B_0_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_522 = _T_43024 ? $signed(_GEN_392) : $signed(TPUs_0_out_B_0_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_523 = _T_43024 ? $signed(_GEN_393) : $signed(TPUs_0_out_B_0_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_524 = _T_43024 ? $signed(_GEN_394) : $signed(TPUs_0_out_B_1_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_525 = _T_43024 ? $signed(_GEN_395) : $signed(TPUs_0_out_B_1_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_526 = _T_43024 ? $signed(_GEN_396) : $signed(TPUs_0_out_B_1_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_527 = _T_43024 ? $signed(_GEN_397) : $signed(TPUs_0_out_B_1_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_528 = _T_43024 ? $signed(_GEN_398) : $signed(TPUs_0_out_B_1_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_529 = _T_43024 ? $signed(_GEN_399) : $signed(TPUs_0_out_B_1_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_530 = _T_43024 ? $signed(_GEN_400) : $signed(TPUs_0_out_B_1_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_531 = _T_43024 ? $signed(_GEN_401) : $signed(TPUs_0_out_B_1_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_532 = _T_43024 ? $signed(_GEN_402) : $signed(TPUs_0_out_B_2_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_533 = _T_43024 ? $signed(_GEN_403) : $signed(TPUs_0_out_B_2_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_534 = _T_43024 ? $signed(_GEN_404) : $signed(TPUs_0_out_B_2_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_535 = _T_43024 ? $signed(_GEN_405) : $signed(TPUs_0_out_B_2_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_536 = _T_43024 ? $signed(_GEN_406) : $signed(TPUs_0_out_B_2_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_537 = _T_43024 ? $signed(_GEN_407) : $signed(TPUs_0_out_B_2_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_538 = _T_43024 ? $signed(_GEN_408) : $signed(TPUs_0_out_B_2_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_539 = _T_43024 ? $signed(_GEN_409) : $signed(TPUs_0_out_B_2_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_540 = _T_43024 ? $signed(_GEN_410) : $signed(TPUs_0_out_B_3_0); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_541 = _T_43024 ? $signed(_GEN_411) : $signed(TPUs_0_out_B_3_1); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_542 = _T_43024 ? $signed(_GEN_412) : $signed(TPUs_0_out_B_3_2); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_543 = _T_43024 ? $signed(_GEN_413) : $signed(TPUs_0_out_B_3_3); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_544 = _T_43024 ? $signed(_GEN_414) : $signed(TPUs_0_out_B_3_4); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_545 = _T_43024 ? $signed(_GEN_415) : $signed(TPUs_0_out_B_3_5); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_546 = _T_43024 ? $signed(_GEN_416) : $signed(TPUs_0_out_B_3_6); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_547 = _T_43024 ? $signed(_GEN_417) : $signed(TPUs_0_out_B_3_7); // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_580 = _T_43024 ? _GEN_208 : TPUs_0_out_tag_0_0; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_581 = _T_43024 ? _GEN_209 : TPUs_0_out_tag_0_1; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_582 = _T_43024 ? _GEN_210 : TPUs_0_out_tag_0_2; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_583 = _T_43024 ? _GEN_211 : TPUs_0_out_tag_0_3; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_584 = _T_43024 ? _GEN_212 : TPUs_0_out_tag_0_4; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_585 = _T_43024 ? _GEN_213 : TPUs_0_out_tag_0_5; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_586 = _T_43024 ? _GEN_214 : TPUs_0_out_tag_0_6; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_587 = _T_43024 ? _GEN_215 : TPUs_0_out_tag_0_7; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_588 = _T_43024 ? _GEN_216 : TPUs_0_out_tag_1_0; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_589 = _T_43024 ? _GEN_217 : TPUs_0_out_tag_1_1; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_590 = _T_43024 ? _GEN_218 : TPUs_0_out_tag_1_2; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_591 = _T_43024 ? _GEN_219 : TPUs_0_out_tag_1_3; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_592 = _T_43024 ? _GEN_220 : TPUs_0_out_tag_1_4; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_593 = _T_43024 ? _GEN_221 : TPUs_0_out_tag_1_5; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_594 = _T_43024 ? _GEN_222 : TPUs_0_out_tag_1_6; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_595 = _T_43024 ? _GEN_223 : TPUs_0_out_tag_1_7; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_596 = _T_43024 ? _GEN_224 : TPUs_0_out_tag_2_0; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_597 = _T_43024 ? _GEN_225 : TPUs_0_out_tag_2_1; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_598 = _T_43024 ? _GEN_226 : TPUs_0_out_tag_2_2; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_599 = _T_43024 ? _GEN_227 : TPUs_0_out_tag_2_3; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_600 = _T_43024 ? _GEN_228 : TPUs_0_out_tag_2_4; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_601 = _T_43024 ? _GEN_229 : TPUs_0_out_tag_2_5; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_602 = _T_43024 ? _GEN_230 : TPUs_0_out_tag_2_6; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_603 = _T_43024 ? _GEN_231 : TPUs_0_out_tag_2_7; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_604 = _T_43024 ? _GEN_232 : TPUs_0_out_tag_3_0; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_605 = _T_43024 ? _GEN_233 : TPUs_0_out_tag_3_1; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_606 = _T_43024 ? _GEN_234 : TPUs_0_out_tag_3_2; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_607 = _T_43024 ? _GEN_235 : TPUs_0_out_tag_3_3; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_608 = _T_43024 ? _GEN_236 : TPUs_0_out_tag_3_4; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_609 = _T_43024 ? _GEN_237 : TPUs_0_out_tag_3_5; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_610 = _T_43024 ? _GEN_238 : TPUs_0_out_tag_3_6; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_611 = _T_43024 ? _GEN_239 : TPUs_0_out_tag_3_7; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_612 = _T_43024 ? _GEN_240 : _GEN_496; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_613 = _T_43024 ? _GEN_241 : cal_control_1; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_614 = _T_43024 ? _GEN_484 : _GEN_499; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_615 = _T_43024 ? cal_control_2 : _GEN_497; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_616 = _T_43024 ? cal_control_0 : _GEN_498; // @[Conditional.scala 39:67:@10413.12]
  assign _GEN_617 = _T_43016 ? $signed(_GEN_250) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_618 = _T_43016 ? $signed(_GEN_251) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_619 = _T_43016 ? $signed(_GEN_252) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_620 = _T_43016 ? $signed(_GEN_253) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_621 = _T_43016 ? $signed(_GEN_254) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_622 = _T_43016 ? $signed(_GEN_255) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_623 = _T_43016 ? $signed(_GEN_256) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_624 = _T_43016 ? $signed(_GEN_257) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_625 = _T_43016 ? $signed(_GEN_258) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_626 = _T_43016 ? $signed(_GEN_259) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_627 = _T_43016 ? $signed(_GEN_260) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_628 = _T_43016 ? $signed(_GEN_261) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_629 = _T_43016 ? $signed(_GEN_262) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_630 = _T_43016 ? $signed(_GEN_263) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_631 = _T_43016 ? $signed(_GEN_264) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_632 = _T_43016 ? $signed(_GEN_265) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_633 = _T_43016 ? $signed(_GEN_266) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_634 = _T_43016 ? $signed(_GEN_267) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_635 = _T_43016 ? $signed(_GEN_268) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_636 = _T_43016 ? $signed(_GEN_269) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_637 = _T_43016 ? $signed(_GEN_270) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_638 = _T_43016 ? $signed(_GEN_271) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_639 = _T_43016 ? $signed(_GEN_272) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_640 = _T_43016 ? $signed(_GEN_273) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_641 = _T_43016 ? $signed(_GEN_274) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_642 = _T_43016 ? $signed(_GEN_275) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_643 = _T_43016 ? $signed(_GEN_276) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_644 = _T_43016 ? $signed(_GEN_277) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_645 = _T_43016 ? $signed(_GEN_278) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_646 = _T_43016 ? $signed(_GEN_279) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_647 = _T_43016 ? $signed(_GEN_280) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_648 = _T_43016 ? $signed(_GEN_281) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_649 = _T_43016 ? $signed(_GEN_282) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_650 = _T_43016 ? $signed(_GEN_283) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_651 = _T_43016 ? $signed(_GEN_284) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_652 = _T_43016 ? $signed(_GEN_285) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_653 = _T_43016 ? $signed(_GEN_286) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_654 = _T_43016 ? $signed(_GEN_287) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_655 = _T_43016 ? $signed(_GEN_288) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_656 = _T_43016 ? $signed(_GEN_289) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_657 = _T_43016 ? $signed(_GEN_290) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_658 = _T_43016 ? $signed(_GEN_291) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_659 = _T_43016 ? $signed(_GEN_292) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_660 = _T_43016 ? $signed(_GEN_293) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_661 = _T_43016 ? $signed(_GEN_294) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_662 = _T_43016 ? $signed(_GEN_295) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_663 = _T_43016 ? $signed(_GEN_296) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_664 = _T_43016 ? $signed(_GEN_297) : $signed(32'sh0); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_729 = _T_43016 ? _GEN_362 : _GEN_612; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_730 = _T_43016 ? _GEN_363 : _GEN_616; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_731 = _T_43016 ? _GEN_364 : _GEN_615; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_732 = _T_43016 ? _GEN_365 : _GEN_614; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_733 = _T_43016 ? $signed(TPUs_0_out_A_0_0) : $signed(_GEN_500); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_734 = _T_43016 ? $signed(TPUs_0_out_A_0_1) : $signed(_GEN_501); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_735 = _T_43016 ? $signed(TPUs_0_out_A_0_2) : $signed(_GEN_502); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_736 = _T_43016 ? $signed(TPUs_0_out_A_0_3) : $signed(_GEN_503); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_737 = _T_43016 ? $signed(TPUs_0_out_A_0_4) : $signed(_GEN_504); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_738 = _T_43016 ? $signed(TPUs_0_out_A_0_5) : $signed(_GEN_505); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_739 = _T_43016 ? $signed(TPUs_0_out_A_0_6) : $signed(_GEN_506); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_740 = _T_43016 ? $signed(TPUs_0_out_A_0_7) : $signed(_GEN_507); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_741 = _T_43016 ? $signed(TPUs_0_out_A_1_0) : $signed(_GEN_508); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_742 = _T_43016 ? $signed(TPUs_0_out_A_1_1) : $signed(_GEN_509); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_743 = _T_43016 ? $signed(TPUs_0_out_A_1_2) : $signed(_GEN_510); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_744 = _T_43016 ? $signed(TPUs_0_out_A_1_3) : $signed(_GEN_511); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_745 = _T_43016 ? $signed(TPUs_0_out_A_1_4) : $signed(_GEN_512); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_746 = _T_43016 ? $signed(TPUs_0_out_A_1_5) : $signed(_GEN_513); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_747 = _T_43016 ? $signed(TPUs_0_out_A_1_6) : $signed(_GEN_514); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_748 = _T_43016 ? $signed(TPUs_0_out_A_1_7) : $signed(_GEN_515); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_749 = _T_43016 ? $signed(TPUs_0_out_B_0_0) : $signed(_GEN_516); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_750 = _T_43016 ? $signed(TPUs_0_out_B_0_1) : $signed(_GEN_517); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_751 = _T_43016 ? $signed(TPUs_0_out_B_0_2) : $signed(_GEN_518); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_752 = _T_43016 ? $signed(TPUs_0_out_B_0_3) : $signed(_GEN_519); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_753 = _T_43016 ? $signed(TPUs_0_out_B_0_4) : $signed(_GEN_520); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_754 = _T_43016 ? $signed(TPUs_0_out_B_0_5) : $signed(_GEN_521); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_755 = _T_43016 ? $signed(TPUs_0_out_B_0_6) : $signed(_GEN_522); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_756 = _T_43016 ? $signed(TPUs_0_out_B_0_7) : $signed(_GEN_523); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_757 = _T_43016 ? $signed(TPUs_0_out_B_1_0) : $signed(_GEN_524); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_758 = _T_43016 ? $signed(TPUs_0_out_B_1_1) : $signed(_GEN_525); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_759 = _T_43016 ? $signed(TPUs_0_out_B_1_2) : $signed(_GEN_526); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_760 = _T_43016 ? $signed(TPUs_0_out_B_1_3) : $signed(_GEN_527); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_761 = _T_43016 ? $signed(TPUs_0_out_B_1_4) : $signed(_GEN_528); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_762 = _T_43016 ? $signed(TPUs_0_out_B_1_5) : $signed(_GEN_529); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_763 = _T_43016 ? $signed(TPUs_0_out_B_1_6) : $signed(_GEN_530); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_764 = _T_43016 ? $signed(TPUs_0_out_B_1_7) : $signed(_GEN_531); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_765 = _T_43016 ? $signed(TPUs_0_out_B_2_0) : $signed(_GEN_532); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_766 = _T_43016 ? $signed(TPUs_0_out_B_2_1) : $signed(_GEN_533); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_767 = _T_43016 ? $signed(TPUs_0_out_B_2_2) : $signed(_GEN_534); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_768 = _T_43016 ? $signed(TPUs_0_out_B_2_3) : $signed(_GEN_535); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_769 = _T_43016 ? $signed(TPUs_0_out_B_2_4) : $signed(_GEN_536); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_770 = _T_43016 ? $signed(TPUs_0_out_B_2_5) : $signed(_GEN_537); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_771 = _T_43016 ? $signed(TPUs_0_out_B_2_6) : $signed(_GEN_538); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_772 = _T_43016 ? $signed(TPUs_0_out_B_2_7) : $signed(_GEN_539); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_773 = _T_43016 ? $signed(TPUs_0_out_B_3_0) : $signed(_GEN_540); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_774 = _T_43016 ? $signed(TPUs_0_out_B_3_1) : $signed(_GEN_541); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_775 = _T_43016 ? $signed(TPUs_0_out_B_3_2) : $signed(_GEN_542); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_776 = _T_43016 ? $signed(TPUs_0_out_B_3_3) : $signed(_GEN_543); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_777 = _T_43016 ? $signed(TPUs_0_out_B_3_4) : $signed(_GEN_544); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_778 = _T_43016 ? $signed(TPUs_0_out_B_3_5) : $signed(_GEN_545); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_779 = _T_43016 ? $signed(TPUs_0_out_B_3_6) : $signed(_GEN_546); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_780 = _T_43016 ? $signed(TPUs_0_out_B_3_7) : $signed(_GEN_547); // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_781 = _T_43016 ? TPUs_0_out_tag_0_0 : _GEN_580; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_782 = _T_43016 ? TPUs_0_out_tag_0_1 : _GEN_581; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_783 = _T_43016 ? TPUs_0_out_tag_0_2 : _GEN_582; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_784 = _T_43016 ? TPUs_0_out_tag_0_3 : _GEN_583; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_785 = _T_43016 ? TPUs_0_out_tag_0_4 : _GEN_584; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_786 = _T_43016 ? TPUs_0_out_tag_0_5 : _GEN_585; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_787 = _T_43016 ? TPUs_0_out_tag_0_6 : _GEN_586; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_788 = _T_43016 ? TPUs_0_out_tag_0_7 : _GEN_587; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_789 = _T_43016 ? TPUs_0_out_tag_1_0 : _GEN_588; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_790 = _T_43016 ? TPUs_0_out_tag_1_1 : _GEN_589; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_791 = _T_43016 ? TPUs_0_out_tag_1_2 : _GEN_590; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_792 = _T_43016 ? TPUs_0_out_tag_1_3 : _GEN_591; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_793 = _T_43016 ? TPUs_0_out_tag_1_4 : _GEN_592; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_794 = _T_43016 ? TPUs_0_out_tag_1_5 : _GEN_593; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_795 = _T_43016 ? TPUs_0_out_tag_1_6 : _GEN_594; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_796 = _T_43016 ? TPUs_0_out_tag_1_7 : _GEN_595; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_797 = _T_43016 ? TPUs_0_out_tag_2_0 : _GEN_596; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_798 = _T_43016 ? TPUs_0_out_tag_2_1 : _GEN_597; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_799 = _T_43016 ? TPUs_0_out_tag_2_2 : _GEN_598; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_800 = _T_43016 ? TPUs_0_out_tag_2_3 : _GEN_599; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_801 = _T_43016 ? TPUs_0_out_tag_2_4 : _GEN_600; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_802 = _T_43016 ? TPUs_0_out_tag_2_5 : _GEN_601; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_803 = _T_43016 ? TPUs_0_out_tag_2_6 : _GEN_602; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_804 = _T_43016 ? TPUs_0_out_tag_2_7 : _GEN_603; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_805 = _T_43016 ? TPUs_0_out_tag_3_0 : _GEN_604; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_806 = _T_43016 ? TPUs_0_out_tag_3_1 : _GEN_605; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_807 = _T_43016 ? TPUs_0_out_tag_3_2 : _GEN_606; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_808 = _T_43016 ? TPUs_0_out_tag_3_3 : _GEN_607; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_809 = _T_43016 ? TPUs_0_out_tag_3_4 : _GEN_608; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_810 = _T_43016 ? TPUs_0_out_tag_3_5 : _GEN_609; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_811 = _T_43016 ? TPUs_0_out_tag_3_6 : _GEN_610; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_812 = _T_43016 ? TPUs_0_out_tag_3_7 : _GEN_611; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_813 = _T_43016 ? cal_control_1 : _GEN_613; // @[Conditional.scala 39:67:@10280.10]
  assign _GEN_814 = _T_43011 ? $signed(_GEN_128) : $signed(_GEN_733); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_815 = _T_43011 ? $signed(_GEN_129) : $signed(_GEN_734); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_816 = _T_43011 ? $signed(_GEN_130) : $signed(_GEN_735); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_817 = _T_43011 ? $signed(_GEN_131) : $signed(_GEN_736); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_818 = _T_43011 ? $signed(_GEN_132) : $signed(_GEN_737); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_819 = _T_43011 ? $signed(_GEN_133) : $signed(_GEN_738); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_820 = _T_43011 ? $signed(_GEN_134) : $signed(_GEN_739); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_821 = _T_43011 ? $signed(_GEN_135) : $signed(_GEN_740); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_822 = _T_43011 ? $signed(_GEN_136) : $signed(_GEN_741); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_823 = _T_43011 ? $signed(_GEN_137) : $signed(_GEN_742); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_824 = _T_43011 ? $signed(_GEN_138) : $signed(_GEN_743); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_825 = _T_43011 ? $signed(_GEN_139) : $signed(_GEN_744); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_826 = _T_43011 ? $signed(_GEN_140) : $signed(_GEN_745); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_827 = _T_43011 ? $signed(_GEN_141) : $signed(_GEN_746); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_828 = _T_43011 ? $signed(_GEN_142) : $signed(_GEN_747); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_829 = _T_43011 ? $signed(_GEN_143) : $signed(_GEN_748); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_830 = _T_43011 ? $signed(_GEN_144) : $signed(_GEN_749); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_831 = _T_43011 ? $signed(_GEN_145) : $signed(_GEN_750); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_832 = _T_43011 ? $signed(_GEN_146) : $signed(_GEN_751); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_833 = _T_43011 ? $signed(_GEN_147) : $signed(_GEN_752); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_834 = _T_43011 ? $signed(_GEN_148) : $signed(_GEN_753); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_835 = _T_43011 ? $signed(_GEN_149) : $signed(_GEN_754); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_836 = _T_43011 ? $signed(_GEN_150) : $signed(_GEN_755); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_837 = _T_43011 ? $signed(_GEN_151) : $signed(_GEN_756); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_838 = _T_43011 ? $signed(_GEN_152) : $signed(_GEN_757); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_839 = _T_43011 ? $signed(_GEN_153) : $signed(_GEN_758); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_840 = _T_43011 ? $signed(_GEN_154) : $signed(_GEN_759); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_841 = _T_43011 ? $signed(_GEN_155) : $signed(_GEN_760); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_842 = _T_43011 ? $signed(_GEN_156) : $signed(_GEN_761); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_843 = _T_43011 ? $signed(_GEN_157) : $signed(_GEN_762); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_844 = _T_43011 ? $signed(_GEN_158) : $signed(_GEN_763); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_845 = _T_43011 ? $signed(_GEN_159) : $signed(_GEN_764); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_846 = _T_43011 ? $signed(_GEN_160) : $signed(_GEN_765); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_847 = _T_43011 ? $signed(_GEN_161) : $signed(_GEN_766); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_848 = _T_43011 ? $signed(_GEN_162) : $signed(_GEN_767); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_849 = _T_43011 ? $signed(_GEN_163) : $signed(_GEN_768); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_850 = _T_43011 ? $signed(_GEN_164) : $signed(_GEN_769); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_851 = _T_43011 ? $signed(_GEN_165) : $signed(_GEN_770); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_852 = _T_43011 ? $signed(_GEN_166) : $signed(_GEN_771); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_853 = _T_43011 ? $signed(_GEN_167) : $signed(_GEN_772); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_854 = _T_43011 ? $signed(_GEN_168) : $signed(_GEN_773); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_855 = _T_43011 ? $signed(_GEN_169) : $signed(_GEN_774); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_856 = _T_43011 ? $signed(_GEN_170) : $signed(_GEN_775); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_857 = _T_43011 ? $signed(_GEN_171) : $signed(_GEN_776); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_858 = _T_43011 ? $signed(_GEN_172) : $signed(_GEN_777); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_859 = _T_43011 ? $signed(_GEN_173) : $signed(_GEN_778); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_860 = _T_43011 ? $signed(_GEN_174) : $signed(_GEN_779); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_861 = _T_43011 ? $signed(_GEN_175) : $signed(_GEN_780); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_894 = _T_43011 ? _GEN_208 : _GEN_781; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_895 = _T_43011 ? _GEN_209 : _GEN_782; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_896 = _T_43011 ? _GEN_210 : _GEN_783; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_897 = _T_43011 ? _GEN_211 : _GEN_784; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_898 = _T_43011 ? _GEN_212 : _GEN_785; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_899 = _T_43011 ? _GEN_213 : _GEN_786; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_900 = _T_43011 ? _GEN_214 : _GEN_787; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_901 = _T_43011 ? _GEN_215 : _GEN_788; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_902 = _T_43011 ? _GEN_216 : _GEN_789; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_903 = _T_43011 ? _GEN_217 : _GEN_790; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_904 = _T_43011 ? _GEN_218 : _GEN_791; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_905 = _T_43011 ? _GEN_219 : _GEN_792; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_906 = _T_43011 ? _GEN_220 : _GEN_793; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_907 = _T_43011 ? _GEN_221 : _GEN_794; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_908 = _T_43011 ? _GEN_222 : _GEN_795; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_909 = _T_43011 ? _GEN_223 : _GEN_796; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_910 = _T_43011 ? _GEN_224 : _GEN_797; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_911 = _T_43011 ? _GEN_225 : _GEN_798; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_912 = _T_43011 ? _GEN_226 : _GEN_799; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_913 = _T_43011 ? _GEN_227 : _GEN_800; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_914 = _T_43011 ? _GEN_228 : _GEN_801; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_915 = _T_43011 ? _GEN_229 : _GEN_802; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_916 = _T_43011 ? _GEN_230 : _GEN_803; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_917 = _T_43011 ? _GEN_231 : _GEN_804; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_918 = _T_43011 ? _GEN_232 : _GEN_805; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_919 = _T_43011 ? _GEN_233 : _GEN_806; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_920 = _T_43011 ? _GEN_234 : _GEN_807; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_921 = _T_43011 ? _GEN_235 : _GEN_808; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_922 = _T_43011 ? _GEN_236 : _GEN_809; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_923 = _T_43011 ? _GEN_237 : _GEN_810; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_924 = _T_43011 ? _GEN_238 : _GEN_811; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_925 = _T_43011 ? _GEN_239 : _GEN_812; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_926 = _T_43011 ? _GEN_240 : _GEN_729; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_927 = _T_43011 ? _GEN_241 : _GEN_813; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_928 = _T_43011 ? _GEN_242 : _GEN_732; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_929 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_617); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_930 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_618); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_931 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_619); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_932 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_620); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_933 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_621); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_934 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_622); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_935 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_623); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_936 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_624); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_937 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_625); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_938 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_626); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_939 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_627); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_940 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_628); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_941 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_629); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_942 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_630); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_943 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_631); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_944 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_632); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_945 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_633); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_946 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_634); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_947 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_635); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_948 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_636); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_949 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_637); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_950 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_638); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_951 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_639); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_952 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_640); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_953 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_641); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_954 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_642); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_955 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_643); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_956 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_644); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_957 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_645); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_958 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_646); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_959 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_647); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_960 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_648); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_961 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_649); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_962 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_650); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_963 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_651); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_964 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_652); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_965 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_653); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_966 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_654); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_967 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_655); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_968 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_656); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_969 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_657); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_970 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_658); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_971 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_659); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_972 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_660); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_973 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_661); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_974 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_662); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_975 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_663); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_976 = _T_43011 ? $signed(32'sh0) : $signed(_GEN_664); // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_1009 = _T_43011 ? cal_control_0 : _GEN_730; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_1010 = _T_43011 ? cal_control_2 : _GEN_731; // @[Conditional.scala 39:67:@10150.8]
  assign _GEN_1011 = _T_43006 ? $signed(_GEN_7) : $signed(_GEN_929); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1012 = _T_43006 ? $signed(_GEN_8) : $signed(_GEN_930); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1013 = _T_43006 ? $signed(_GEN_9) : $signed(_GEN_931); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1014 = _T_43006 ? $signed(_GEN_10) : $signed(_GEN_932); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1015 = _T_43006 ? $signed(_GEN_11) : $signed(_GEN_933); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1016 = _T_43006 ? $signed(_GEN_12) : $signed(_GEN_934); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1017 = _T_43006 ? $signed(_GEN_13) : $signed(_GEN_935); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1018 = _T_43006 ? $signed(_GEN_14) : $signed(_GEN_936); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1019 = _T_43006 ? $signed(_GEN_15) : $signed(_GEN_937); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1020 = _T_43006 ? $signed(_GEN_16) : $signed(_GEN_938); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1021 = _T_43006 ? $signed(_GEN_17) : $signed(_GEN_939); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1022 = _T_43006 ? $signed(_GEN_18) : $signed(_GEN_940); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1023 = _T_43006 ? $signed(_GEN_19) : $signed(_GEN_941); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1024 = _T_43006 ? $signed(_GEN_20) : $signed(_GEN_942); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1025 = _T_43006 ? $signed(_GEN_21) : $signed(_GEN_943); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1026 = _T_43006 ? $signed(_GEN_22) : $signed(_GEN_944); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1027 = _T_43006 ? $signed(_GEN_23) : $signed(_GEN_945); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1028 = _T_43006 ? $signed(_GEN_24) : $signed(_GEN_946); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1029 = _T_43006 ? $signed(_GEN_25) : $signed(_GEN_947); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1030 = _T_43006 ? $signed(_GEN_26) : $signed(_GEN_948); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1031 = _T_43006 ? $signed(_GEN_27) : $signed(_GEN_949); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1032 = _T_43006 ? $signed(_GEN_28) : $signed(_GEN_950); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1033 = _T_43006 ? $signed(_GEN_29) : $signed(_GEN_951); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1034 = _T_43006 ? $signed(_GEN_30) : $signed(_GEN_952); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1035 = _T_43006 ? $signed(_GEN_31) : $signed(_GEN_953); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1036 = _T_43006 ? $signed(_GEN_32) : $signed(_GEN_954); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1037 = _T_43006 ? $signed(_GEN_33) : $signed(_GEN_955); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1038 = _T_43006 ? $signed(_GEN_34) : $signed(_GEN_956); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1039 = _T_43006 ? $signed(_GEN_35) : $signed(_GEN_957); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1040 = _T_43006 ? $signed(_GEN_36) : $signed(_GEN_958); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1041 = _T_43006 ? $signed(_GEN_37) : $signed(_GEN_959); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1042 = _T_43006 ? $signed(_GEN_38) : $signed(_GEN_960); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1043 = _T_43006 ? $signed(_GEN_39) : $signed(_GEN_961); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1044 = _T_43006 ? $signed(_GEN_40) : $signed(_GEN_962); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1045 = _T_43006 ? $signed(_GEN_41) : $signed(_GEN_963); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1046 = _T_43006 ? $signed(_GEN_42) : $signed(_GEN_964); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1047 = _T_43006 ? $signed(_GEN_43) : $signed(_GEN_965); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1048 = _T_43006 ? $signed(_GEN_44) : $signed(_GEN_966); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1049 = _T_43006 ? $signed(_GEN_45) : $signed(_GEN_967); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1050 = _T_43006 ? $signed(_GEN_46) : $signed(_GEN_968); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1051 = _T_43006 ? $signed(_GEN_47) : $signed(_GEN_969); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1052 = _T_43006 ? $signed(_GEN_48) : $signed(_GEN_970); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1053 = _T_43006 ? $signed(_GEN_49) : $signed(_GEN_971); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1054 = _T_43006 ? $signed(_GEN_50) : $signed(_GEN_972); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1055 = _T_43006 ? $signed(_GEN_51) : $signed(_GEN_973); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1056 = _T_43006 ? $signed(_GEN_52) : $signed(_GEN_974); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1057 = _T_43006 ? $signed(_GEN_53) : $signed(_GEN_975); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1058 = _T_43006 ? $signed(_GEN_54) : $signed(_GEN_976); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1123 = _T_43006 ? _GEN_119 : _GEN_926; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1124 = _T_43006 ? _GEN_120 : _GEN_1009; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1125 = _T_43006 ? _GEN_121 : _GEN_928; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1126 = _T_43006 ? $signed(TPUs_0_out_A_0_0) : $signed(_GEN_814); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1127 = _T_43006 ? $signed(TPUs_0_out_A_0_1) : $signed(_GEN_815); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1128 = _T_43006 ? $signed(TPUs_0_out_A_0_2) : $signed(_GEN_816); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1129 = _T_43006 ? $signed(TPUs_0_out_A_0_3) : $signed(_GEN_817); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1130 = _T_43006 ? $signed(TPUs_0_out_A_0_4) : $signed(_GEN_818); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1131 = _T_43006 ? $signed(TPUs_0_out_A_0_5) : $signed(_GEN_819); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1132 = _T_43006 ? $signed(TPUs_0_out_A_0_6) : $signed(_GEN_820); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1133 = _T_43006 ? $signed(TPUs_0_out_A_0_7) : $signed(_GEN_821); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1134 = _T_43006 ? $signed(TPUs_0_out_A_1_0) : $signed(_GEN_822); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1135 = _T_43006 ? $signed(TPUs_0_out_A_1_1) : $signed(_GEN_823); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1136 = _T_43006 ? $signed(TPUs_0_out_A_1_2) : $signed(_GEN_824); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1137 = _T_43006 ? $signed(TPUs_0_out_A_1_3) : $signed(_GEN_825); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1138 = _T_43006 ? $signed(TPUs_0_out_A_1_4) : $signed(_GEN_826); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1139 = _T_43006 ? $signed(TPUs_0_out_A_1_5) : $signed(_GEN_827); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1140 = _T_43006 ? $signed(TPUs_0_out_A_1_6) : $signed(_GEN_828); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1141 = _T_43006 ? $signed(TPUs_0_out_A_1_7) : $signed(_GEN_829); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1142 = _T_43006 ? $signed(TPUs_0_out_B_0_0) : $signed(_GEN_830); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1143 = _T_43006 ? $signed(TPUs_0_out_B_0_1) : $signed(_GEN_831); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1144 = _T_43006 ? $signed(TPUs_0_out_B_0_2) : $signed(_GEN_832); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1145 = _T_43006 ? $signed(TPUs_0_out_B_0_3) : $signed(_GEN_833); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1146 = _T_43006 ? $signed(TPUs_0_out_B_0_4) : $signed(_GEN_834); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1147 = _T_43006 ? $signed(TPUs_0_out_B_0_5) : $signed(_GEN_835); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1148 = _T_43006 ? $signed(TPUs_0_out_B_0_6) : $signed(_GEN_836); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1149 = _T_43006 ? $signed(TPUs_0_out_B_0_7) : $signed(_GEN_837); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1150 = _T_43006 ? $signed(TPUs_0_out_B_1_0) : $signed(_GEN_838); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1151 = _T_43006 ? $signed(TPUs_0_out_B_1_1) : $signed(_GEN_839); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1152 = _T_43006 ? $signed(TPUs_0_out_B_1_2) : $signed(_GEN_840); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1153 = _T_43006 ? $signed(TPUs_0_out_B_1_3) : $signed(_GEN_841); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1154 = _T_43006 ? $signed(TPUs_0_out_B_1_4) : $signed(_GEN_842); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1155 = _T_43006 ? $signed(TPUs_0_out_B_1_5) : $signed(_GEN_843); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1156 = _T_43006 ? $signed(TPUs_0_out_B_1_6) : $signed(_GEN_844); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1157 = _T_43006 ? $signed(TPUs_0_out_B_1_7) : $signed(_GEN_845); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1158 = _T_43006 ? $signed(TPUs_0_out_B_2_0) : $signed(_GEN_846); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1159 = _T_43006 ? $signed(TPUs_0_out_B_2_1) : $signed(_GEN_847); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1160 = _T_43006 ? $signed(TPUs_0_out_B_2_2) : $signed(_GEN_848); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1161 = _T_43006 ? $signed(TPUs_0_out_B_2_3) : $signed(_GEN_849); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1162 = _T_43006 ? $signed(TPUs_0_out_B_2_4) : $signed(_GEN_850); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1163 = _T_43006 ? $signed(TPUs_0_out_B_2_5) : $signed(_GEN_851); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1164 = _T_43006 ? $signed(TPUs_0_out_B_2_6) : $signed(_GEN_852); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1165 = _T_43006 ? $signed(TPUs_0_out_B_2_7) : $signed(_GEN_853); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1166 = _T_43006 ? $signed(TPUs_0_out_B_3_0) : $signed(_GEN_854); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1167 = _T_43006 ? $signed(TPUs_0_out_B_3_1) : $signed(_GEN_855); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1168 = _T_43006 ? $signed(TPUs_0_out_B_3_2) : $signed(_GEN_856); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1169 = _T_43006 ? $signed(TPUs_0_out_B_3_3) : $signed(_GEN_857); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1170 = _T_43006 ? $signed(TPUs_0_out_B_3_4) : $signed(_GEN_858); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1171 = _T_43006 ? $signed(TPUs_0_out_B_3_5) : $signed(_GEN_859); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1172 = _T_43006 ? $signed(TPUs_0_out_B_3_6) : $signed(_GEN_860); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1173 = _T_43006 ? $signed(TPUs_0_out_B_3_7) : $signed(_GEN_861); // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1174 = _T_43006 ? TPUs_0_out_tag_0_0 : _GEN_894; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1175 = _T_43006 ? TPUs_0_out_tag_0_1 : _GEN_895; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1176 = _T_43006 ? TPUs_0_out_tag_0_2 : _GEN_896; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1177 = _T_43006 ? TPUs_0_out_tag_0_3 : _GEN_897; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1178 = _T_43006 ? TPUs_0_out_tag_0_4 : _GEN_898; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1179 = _T_43006 ? TPUs_0_out_tag_0_5 : _GEN_899; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1180 = _T_43006 ? TPUs_0_out_tag_0_6 : _GEN_900; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1181 = _T_43006 ? TPUs_0_out_tag_0_7 : _GEN_901; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1182 = _T_43006 ? TPUs_0_out_tag_1_0 : _GEN_902; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1183 = _T_43006 ? TPUs_0_out_tag_1_1 : _GEN_903; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1184 = _T_43006 ? TPUs_0_out_tag_1_2 : _GEN_904; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1185 = _T_43006 ? TPUs_0_out_tag_1_3 : _GEN_905; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1186 = _T_43006 ? TPUs_0_out_tag_1_4 : _GEN_906; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1187 = _T_43006 ? TPUs_0_out_tag_1_5 : _GEN_907; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1188 = _T_43006 ? TPUs_0_out_tag_1_6 : _GEN_908; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1189 = _T_43006 ? TPUs_0_out_tag_1_7 : _GEN_909; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1190 = _T_43006 ? TPUs_0_out_tag_2_0 : _GEN_910; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1191 = _T_43006 ? TPUs_0_out_tag_2_1 : _GEN_911; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1192 = _T_43006 ? TPUs_0_out_tag_2_2 : _GEN_912; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1193 = _T_43006 ? TPUs_0_out_tag_2_3 : _GEN_913; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1194 = _T_43006 ? TPUs_0_out_tag_2_4 : _GEN_914; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1195 = _T_43006 ? TPUs_0_out_tag_2_5 : _GEN_915; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1196 = _T_43006 ? TPUs_0_out_tag_2_6 : _GEN_916; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1197 = _T_43006 ? TPUs_0_out_tag_2_7 : _GEN_917; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1198 = _T_43006 ? TPUs_0_out_tag_3_0 : _GEN_918; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1199 = _T_43006 ? TPUs_0_out_tag_3_1 : _GEN_919; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1200 = _T_43006 ? TPUs_0_out_tag_3_2 : _GEN_920; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1201 = _T_43006 ? TPUs_0_out_tag_3_3 : _GEN_921; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1202 = _T_43006 ? TPUs_0_out_tag_3_4 : _GEN_922; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1203 = _T_43006 ? TPUs_0_out_tag_3_5 : _GEN_923; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1204 = _T_43006 ? TPUs_0_out_tag_3_6 : _GEN_924; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1205 = _T_43006 ? TPUs_0_out_tag_3_7 : _GEN_925; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1206 = _T_43006 ? cal_control_1 : _GEN_927; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1207 = _T_43006 ? cal_control_2 : _GEN_1010; // @[Conditional.scala 39:67:@10020.6]
  assign _GEN_1208 = _T_43000 ? _GEN_0 : _GEN_1125; // @[Conditional.scala 40:58:@10009.4]
  assign _GEN_1321 = _T_43000 ? loop_reg : _GEN_1123; // @[Conditional.scala 40:58:@10009.4]
  assign _GEN_1322 = _T_43000 ? cal_control_0 : _GEN_1124; // @[Conditional.scala 40:58:@10009.4]
  assign _GEN_1403 = _T_43000 ? cal_control_1 : _GEN_1206; // @[Conditional.scala 40:58:@10009.4]
  assign _GEN_1404 = _T_43000 ? cal_control_2 : _GEN_1207; // @[Conditional.scala 40:58:@10009.4]
  assign TPUs_0_out_result_0_0 = TPU_io_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8688.4]
  assign TPUs_0_out_result_0_1 = TPU_io_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8689.4]
  assign TPUs_0_out_result_0_2 = TPU_io_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8690.4]
  assign TPUs_0_out_result_0_3 = TPU_io_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8691.4]
  assign TPUs_0_out_result_1_0 = TPU_io_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8692.4]
  assign TPUs_0_out_result_1_1 = TPU_io_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8693.4]
  assign TPUs_0_out_result_1_2 = TPU_io_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8694.4]
  assign TPUs_0_out_result_1_3 = TPU_io_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8695.4]
  assign TPUs_0_out_cal = TPU_io_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8687.4]
  assign TPUs_1_out_result_0_0 = TPU_1_io_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8858.4]
  assign TPUs_1_out_result_0_1 = TPU_1_io_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8859.4]
  assign TPUs_1_out_result_0_2 = TPU_1_io_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8860.4]
  assign TPUs_1_out_result_0_3 = TPU_1_io_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8861.4]
  assign TPUs_1_out_result_1_0 = TPU_1_io_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8862.4]
  assign TPUs_1_out_result_1_1 = TPU_1_io_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8863.4]
  assign TPUs_1_out_result_1_2 = TPU_1_io_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8864.4]
  assign TPUs_1_out_result_1_3 = TPU_1_io_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@8865.4]
  assign TPUs_2_out_result_0_0 = TPU_2_io_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9028.4]
  assign TPUs_2_out_result_0_1 = TPU_2_io_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9029.4]
  assign TPUs_2_out_result_0_2 = TPU_2_io_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9030.4]
  assign TPUs_2_out_result_0_3 = TPU_2_io_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9031.4]
  assign TPUs_2_out_result_1_0 = TPU_2_io_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9032.4]
  assign TPUs_2_out_result_1_1 = TPU_2_io_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9033.4]
  assign TPUs_2_out_result_1_2 = TPU_2_io_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9034.4]
  assign TPUs_2_out_result_1_3 = TPU_2_io_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9035.4]
  assign TPUs_3_out_result_0_0 = TPU_3_io_out_result_0_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9198.4]
  assign TPUs_3_out_result_0_1 = TPU_3_io_out_result_0_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9199.4]
  assign TPUs_3_out_result_0_2 = TPU_3_io_out_result_0_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9200.4]
  assign TPUs_3_out_result_0_3 = TPU_3_io_out_result_0_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9201.4]
  assign TPUs_3_out_result_1_0 = TPU_3_io_out_result_1_0; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9202.4]
  assign TPUs_3_out_result_1_1 = TPU_3_io_out_result_1_1; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9203.4]
  assign TPUs_3_out_result_1_2 = TPU_3_io_out_result_1_2; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9204.4]
  assign TPUs_3_out_result_1_3 = TPU_3_io_out_result_1_3; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9205.4]
  assign TPUs_3_out_cal = TPU_3_io_out_cal; // @[STA_VDBB.scala 97:17:@8686.4 STA_VDBB.scala 97:17:@9197.4]
  assign io_out_C_0_0 = result_0_0; // @[STA_VDBB.scala 120:12:@9933.4]
  assign io_out_C_0_1 = result_0_1; // @[STA_VDBB.scala 120:12:@9934.4]
  assign io_out_C_0_2 = result_0_2; // @[STA_VDBB.scala 120:12:@9935.4]
  assign io_out_C_0_3 = result_0_3; // @[STA_VDBB.scala 120:12:@9936.4]
  assign io_out_C_0_4 = result_0_4; // @[STA_VDBB.scala 120:12:@9937.4]
  assign io_out_C_0_5 = result_0_5; // @[STA_VDBB.scala 120:12:@9938.4]
  assign io_out_C_0_6 = result_0_6; // @[STA_VDBB.scala 120:12:@9939.4]
  assign io_out_C_0_7 = result_0_7; // @[STA_VDBB.scala 120:12:@9940.4]
  assign io_out_C_1_0 = result_1_0; // @[STA_VDBB.scala 120:12:@9941.4]
  assign io_out_C_1_1 = result_1_1; // @[STA_VDBB.scala 120:12:@9942.4]
  assign io_out_C_1_2 = result_1_2; // @[STA_VDBB.scala 120:12:@9943.4]
  assign io_out_C_1_3 = result_1_3; // @[STA_VDBB.scala 120:12:@9944.4]
  assign io_out_C_1_4 = result_1_4; // @[STA_VDBB.scala 120:12:@9945.4]
  assign io_out_C_1_5 = result_1_5; // @[STA_VDBB.scala 120:12:@9946.4]
  assign io_out_C_1_6 = result_1_6; // @[STA_VDBB.scala 120:12:@9947.4]
  assign io_out_C_1_7 = result_1_7; // @[STA_VDBB.scala 120:12:@9948.4]
  assign io_out_C_2_0 = result_2_0; // @[STA_VDBB.scala 120:12:@9949.4]
  assign io_out_C_2_1 = result_2_1; // @[STA_VDBB.scala 120:12:@9950.4]
  assign io_out_C_2_2 = result_2_2; // @[STA_VDBB.scala 120:12:@9951.4]
  assign io_out_C_2_3 = result_2_3; // @[STA_VDBB.scala 120:12:@9952.4]
  assign io_out_C_2_4 = result_2_4; // @[STA_VDBB.scala 120:12:@9953.4]
  assign io_out_C_2_5 = result_2_5; // @[STA_VDBB.scala 120:12:@9954.4]
  assign io_out_C_2_6 = result_2_6; // @[STA_VDBB.scala 120:12:@9955.4]
  assign io_out_C_2_7 = result_2_7; // @[STA_VDBB.scala 120:12:@9956.4]
  assign io_out_C_3_0 = result_3_0; // @[STA_VDBB.scala 120:12:@9957.4]
  assign io_out_C_3_1 = result_3_1; // @[STA_VDBB.scala 120:12:@9958.4]
  assign io_out_C_3_2 = result_3_2; // @[STA_VDBB.scala 120:12:@9959.4]
  assign io_out_C_3_3 = result_3_3; // @[STA_VDBB.scala 120:12:@9960.4]
  assign io_out_C_3_4 = result_3_4; // @[STA_VDBB.scala 120:12:@9961.4]
  assign io_out_C_3_5 = result_3_5; // @[STA_VDBB.scala 120:12:@9962.4]
  assign io_out_C_3_6 = result_3_6; // @[STA_VDBB.scala 120:12:@9963.4]
  assign io_out_C_3_7 = result_3_7; // @[STA_VDBB.scala 120:12:@9964.4]
  assign io_out_cal = _T_40966 & cal_state_2; // @[STA_VDBB.scala 117:14:@9862.4]
  assign TPU_clock = clock; // @[:@8675.4]
  assign TPU_reset = reset; // @[:@8676.4]
  assign TPU_io_in_A_0_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1011); // @[STA_VDBB.scala 97:17:@8841.4]
  assign TPU_io_in_A_0_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1012); // @[STA_VDBB.scala 97:17:@8842.4]
  assign TPU_io_in_A_0_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1013); // @[STA_VDBB.scala 97:17:@8843.4]
  assign TPU_io_in_A_0_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1014); // @[STA_VDBB.scala 97:17:@8844.4]
  assign TPU_io_in_A_0_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1015); // @[STA_VDBB.scala 97:17:@8845.4]
  assign TPU_io_in_A_0_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1016); // @[STA_VDBB.scala 97:17:@8846.4]
  assign TPU_io_in_A_0_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1017); // @[STA_VDBB.scala 97:17:@8847.4]
  assign TPU_io_in_A_0_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1018); // @[STA_VDBB.scala 97:17:@8848.4]
  assign TPU_io_in_A_1_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1019); // @[STA_VDBB.scala 97:17:@8849.4]
  assign TPU_io_in_A_1_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1020); // @[STA_VDBB.scala 97:17:@8850.4]
  assign TPU_io_in_A_1_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1021); // @[STA_VDBB.scala 97:17:@8851.4]
  assign TPU_io_in_A_1_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1022); // @[STA_VDBB.scala 97:17:@8852.4]
  assign TPU_io_in_A_1_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1023); // @[STA_VDBB.scala 97:17:@8853.4]
  assign TPU_io_in_A_1_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1024); // @[STA_VDBB.scala 97:17:@8854.4]
  assign TPU_io_in_A_1_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1025); // @[STA_VDBB.scala 97:17:@8855.4]
  assign TPU_io_in_A_1_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1026); // @[STA_VDBB.scala 97:17:@8856.4]
  assign TPU_io_in_B_0_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1027); // @[STA_VDBB.scala 97:17:@8809.4]
  assign TPU_io_in_B_0_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1028); // @[STA_VDBB.scala 97:17:@8810.4]
  assign TPU_io_in_B_0_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1029); // @[STA_VDBB.scala 97:17:@8811.4]
  assign TPU_io_in_B_0_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1030); // @[STA_VDBB.scala 97:17:@8812.4]
  assign TPU_io_in_B_0_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1031); // @[STA_VDBB.scala 97:17:@8813.4]
  assign TPU_io_in_B_0_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1032); // @[STA_VDBB.scala 97:17:@8814.4]
  assign TPU_io_in_B_0_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1033); // @[STA_VDBB.scala 97:17:@8815.4]
  assign TPU_io_in_B_0_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1034); // @[STA_VDBB.scala 97:17:@8816.4]
  assign TPU_io_in_B_1_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1035); // @[STA_VDBB.scala 97:17:@8817.4]
  assign TPU_io_in_B_1_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1036); // @[STA_VDBB.scala 97:17:@8818.4]
  assign TPU_io_in_B_1_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1037); // @[STA_VDBB.scala 97:17:@8819.4]
  assign TPU_io_in_B_1_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1038); // @[STA_VDBB.scala 97:17:@8820.4]
  assign TPU_io_in_B_1_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1039); // @[STA_VDBB.scala 97:17:@8821.4]
  assign TPU_io_in_B_1_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1040); // @[STA_VDBB.scala 97:17:@8822.4]
  assign TPU_io_in_B_1_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1041); // @[STA_VDBB.scala 97:17:@8823.4]
  assign TPU_io_in_B_1_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1042); // @[STA_VDBB.scala 97:17:@8824.4]
  assign TPU_io_in_B_2_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1043); // @[STA_VDBB.scala 97:17:@8825.4]
  assign TPU_io_in_B_2_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1044); // @[STA_VDBB.scala 97:17:@8826.4]
  assign TPU_io_in_B_2_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1045); // @[STA_VDBB.scala 97:17:@8827.4]
  assign TPU_io_in_B_2_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1046); // @[STA_VDBB.scala 97:17:@8828.4]
  assign TPU_io_in_B_2_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1047); // @[STA_VDBB.scala 97:17:@8829.4]
  assign TPU_io_in_B_2_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1048); // @[STA_VDBB.scala 97:17:@8830.4]
  assign TPU_io_in_B_2_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1049); // @[STA_VDBB.scala 97:17:@8831.4]
  assign TPU_io_in_B_2_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1050); // @[STA_VDBB.scala 97:17:@8832.4]
  assign TPU_io_in_B_3_0 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1051); // @[STA_VDBB.scala 97:17:@8833.4]
  assign TPU_io_in_B_3_1 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1052); // @[STA_VDBB.scala 97:17:@8834.4]
  assign TPU_io_in_B_3_2 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1053); // @[STA_VDBB.scala 97:17:@8835.4]
  assign TPU_io_in_B_3_3 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1054); // @[STA_VDBB.scala 97:17:@8836.4]
  assign TPU_io_in_B_3_4 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1055); // @[STA_VDBB.scala 97:17:@8837.4]
  assign TPU_io_in_B_3_5 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1056); // @[STA_VDBB.scala 97:17:@8838.4]
  assign TPU_io_in_B_3_6 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1057); // @[STA_VDBB.scala 97:17:@8839.4]
  assign TPU_io_in_B_3_7 = _T_43000 ? $signed(32'sh0) : $signed(_GEN_1058); // @[STA_VDBB.scala 97:17:@8840.4]
  assign TPU_io_in_tag_0_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8777.4]
  assign TPU_io_in_tag_0_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8778.4]
  assign TPU_io_in_tag_0_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8779.4]
  assign TPU_io_in_tag_0_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8780.4]
  assign TPU_io_in_tag_0_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8781.4]
  assign TPU_io_in_tag_0_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8782.4]
  assign TPU_io_in_tag_0_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8783.4]
  assign TPU_io_in_tag_0_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8784.4]
  assign TPU_io_in_tag_1_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8785.4]
  assign TPU_io_in_tag_1_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8786.4]
  assign TPU_io_in_tag_1_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8787.4]
  assign TPU_io_in_tag_1_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8788.4]
  assign TPU_io_in_tag_1_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8789.4]
  assign TPU_io_in_tag_1_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8790.4]
  assign TPU_io_in_tag_1_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8791.4]
  assign TPU_io_in_tag_1_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8792.4]
  assign TPU_io_in_tag_2_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8793.4]
  assign TPU_io_in_tag_2_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8794.4]
  assign TPU_io_in_tag_2_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8795.4]
  assign TPU_io_in_tag_2_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8796.4]
  assign TPU_io_in_tag_2_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8797.4]
  assign TPU_io_in_tag_2_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8798.4]
  assign TPU_io_in_tag_2_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8799.4]
  assign TPU_io_in_tag_2_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8800.4]
  assign TPU_io_in_tag_3_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8801.4]
  assign TPU_io_in_tag_3_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8802.4]
  assign TPU_io_in_tag_3_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8803.4]
  assign TPU_io_in_tag_3_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8804.4]
  assign TPU_io_in_tag_3_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8805.4]
  assign TPU_io_in_tag_3_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8806.4]
  assign TPU_io_in_tag_3_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8807.4]
  assign TPU_io_in_tag_3_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8808.4]
  assign TPU_io_in_cal = cal_control_0; // @[STA_VDBB.scala 97:17:@8776.4]
  assign TPU_1_clock = clock; // @[:@8678.4]
  assign TPU_1_reset = reset; // @[:@8679.4]
  assign TPU_1_io_in_A_0_0 = _T_43000 ? $signed(TPUs_0_out_A_0_0) : $signed(_GEN_1126); // @[STA_VDBB.scala 97:17:@9011.4]
  assign TPU_1_io_in_A_0_1 = _T_43000 ? $signed(TPUs_0_out_A_0_1) : $signed(_GEN_1127); // @[STA_VDBB.scala 97:17:@9012.4]
  assign TPU_1_io_in_A_0_2 = _T_43000 ? $signed(TPUs_0_out_A_0_2) : $signed(_GEN_1128); // @[STA_VDBB.scala 97:17:@9013.4]
  assign TPU_1_io_in_A_0_3 = _T_43000 ? $signed(TPUs_0_out_A_0_3) : $signed(_GEN_1129); // @[STA_VDBB.scala 97:17:@9014.4]
  assign TPU_1_io_in_A_0_4 = _T_43000 ? $signed(TPUs_0_out_A_0_4) : $signed(_GEN_1130); // @[STA_VDBB.scala 97:17:@9015.4]
  assign TPU_1_io_in_A_0_5 = _T_43000 ? $signed(TPUs_0_out_A_0_5) : $signed(_GEN_1131); // @[STA_VDBB.scala 97:17:@9016.4]
  assign TPU_1_io_in_A_0_6 = _T_43000 ? $signed(TPUs_0_out_A_0_6) : $signed(_GEN_1132); // @[STA_VDBB.scala 97:17:@9017.4]
  assign TPU_1_io_in_A_0_7 = _T_43000 ? $signed(TPUs_0_out_A_0_7) : $signed(_GEN_1133); // @[STA_VDBB.scala 97:17:@9018.4]
  assign TPU_1_io_in_A_1_0 = _T_43000 ? $signed(TPUs_0_out_A_1_0) : $signed(_GEN_1134); // @[STA_VDBB.scala 97:17:@9019.4]
  assign TPU_1_io_in_A_1_1 = _T_43000 ? $signed(TPUs_0_out_A_1_1) : $signed(_GEN_1135); // @[STA_VDBB.scala 97:17:@9020.4]
  assign TPU_1_io_in_A_1_2 = _T_43000 ? $signed(TPUs_0_out_A_1_2) : $signed(_GEN_1136); // @[STA_VDBB.scala 97:17:@9021.4]
  assign TPU_1_io_in_A_1_3 = _T_43000 ? $signed(TPUs_0_out_A_1_3) : $signed(_GEN_1137); // @[STA_VDBB.scala 97:17:@9022.4]
  assign TPU_1_io_in_A_1_4 = _T_43000 ? $signed(TPUs_0_out_A_1_4) : $signed(_GEN_1138); // @[STA_VDBB.scala 97:17:@9023.4]
  assign TPU_1_io_in_A_1_5 = _T_43000 ? $signed(TPUs_0_out_A_1_5) : $signed(_GEN_1139); // @[STA_VDBB.scala 97:17:@9024.4]
  assign TPU_1_io_in_A_1_6 = _T_43000 ? $signed(TPUs_0_out_A_1_6) : $signed(_GEN_1140); // @[STA_VDBB.scala 97:17:@9025.4]
  assign TPU_1_io_in_A_1_7 = _T_43000 ? $signed(TPUs_0_out_A_1_7) : $signed(_GEN_1141); // @[STA_VDBB.scala 97:17:@9026.4]
  assign TPU_1_io_in_B_0_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@8979.4]
  assign TPU_1_io_in_B_0_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@8980.4]
  assign TPU_1_io_in_B_0_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@8981.4]
  assign TPU_1_io_in_B_0_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@8982.4]
  assign TPU_1_io_in_B_0_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@8983.4]
  assign TPU_1_io_in_B_0_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@8984.4]
  assign TPU_1_io_in_B_0_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@8985.4]
  assign TPU_1_io_in_B_0_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@8986.4]
  assign TPU_1_io_in_B_1_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@8987.4]
  assign TPU_1_io_in_B_1_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@8988.4]
  assign TPU_1_io_in_B_1_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@8989.4]
  assign TPU_1_io_in_B_1_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@8990.4]
  assign TPU_1_io_in_B_1_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@8991.4]
  assign TPU_1_io_in_B_1_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@8992.4]
  assign TPU_1_io_in_B_1_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@8993.4]
  assign TPU_1_io_in_B_1_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@8994.4]
  assign TPU_1_io_in_B_2_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@8995.4]
  assign TPU_1_io_in_B_2_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@8996.4]
  assign TPU_1_io_in_B_2_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@8997.4]
  assign TPU_1_io_in_B_2_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@8998.4]
  assign TPU_1_io_in_B_2_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@8999.4]
  assign TPU_1_io_in_B_2_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@9000.4]
  assign TPU_1_io_in_B_2_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@9001.4]
  assign TPU_1_io_in_B_2_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@9002.4]
  assign TPU_1_io_in_B_3_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@9003.4]
  assign TPU_1_io_in_B_3_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@9004.4]
  assign TPU_1_io_in_B_3_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@9005.4]
  assign TPU_1_io_in_B_3_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@9006.4]
  assign TPU_1_io_in_B_3_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@9007.4]
  assign TPU_1_io_in_B_3_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@9008.4]
  assign TPU_1_io_in_B_3_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@9009.4]
  assign TPU_1_io_in_B_3_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@9010.4]
  assign TPU_1_io_in_tag_0_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8947.4]
  assign TPU_1_io_in_tag_0_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8948.4]
  assign TPU_1_io_in_tag_0_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8949.4]
  assign TPU_1_io_in_tag_0_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8950.4]
  assign TPU_1_io_in_tag_0_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8951.4]
  assign TPU_1_io_in_tag_0_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8952.4]
  assign TPU_1_io_in_tag_0_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8953.4]
  assign TPU_1_io_in_tag_0_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8954.4]
  assign TPU_1_io_in_tag_1_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8955.4]
  assign TPU_1_io_in_tag_1_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8956.4]
  assign TPU_1_io_in_tag_1_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8957.4]
  assign TPU_1_io_in_tag_1_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8958.4]
  assign TPU_1_io_in_tag_1_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8959.4]
  assign TPU_1_io_in_tag_1_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8960.4]
  assign TPU_1_io_in_tag_1_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8961.4]
  assign TPU_1_io_in_tag_1_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8962.4]
  assign TPU_1_io_in_tag_2_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8963.4]
  assign TPU_1_io_in_tag_2_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8964.4]
  assign TPU_1_io_in_tag_2_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8965.4]
  assign TPU_1_io_in_tag_2_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8966.4]
  assign TPU_1_io_in_tag_2_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8967.4]
  assign TPU_1_io_in_tag_2_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8968.4]
  assign TPU_1_io_in_tag_2_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8969.4]
  assign TPU_1_io_in_tag_2_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8970.4]
  assign TPU_1_io_in_tag_3_0 = 1'h0; // @[STA_VDBB.scala 97:17:@8971.4]
  assign TPU_1_io_in_tag_3_1 = 1'h0; // @[STA_VDBB.scala 97:17:@8972.4]
  assign TPU_1_io_in_tag_3_2 = 1'h0; // @[STA_VDBB.scala 97:17:@8973.4]
  assign TPU_1_io_in_tag_3_3 = 1'h0; // @[STA_VDBB.scala 97:17:@8974.4]
  assign TPU_1_io_in_tag_3_4 = 1'h0; // @[STA_VDBB.scala 97:17:@8975.4]
  assign TPU_1_io_in_tag_3_5 = 1'h0; // @[STA_VDBB.scala 97:17:@8976.4]
  assign TPU_1_io_in_tag_3_6 = 1'h0; // @[STA_VDBB.scala 97:17:@8977.4]
  assign TPU_1_io_in_tag_3_7 = 1'h0; // @[STA_VDBB.scala 97:17:@8978.4]
  assign TPU_1_io_in_cal = cal_control_1; // @[STA_VDBB.scala 97:17:@8946.4]
  assign TPU_2_clock = clock; // @[:@8681.4]
  assign TPU_2_reset = reset; // @[:@8682.4]
  assign TPU_2_io_in_A_0_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@9181.4]
  assign TPU_2_io_in_A_0_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@9182.4]
  assign TPU_2_io_in_A_0_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@9183.4]
  assign TPU_2_io_in_A_0_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@9184.4]
  assign TPU_2_io_in_A_0_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@9185.4]
  assign TPU_2_io_in_A_0_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@9186.4]
  assign TPU_2_io_in_A_0_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@9187.4]
  assign TPU_2_io_in_A_0_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@9188.4]
  assign TPU_2_io_in_A_1_0 = 32'sh0; // @[STA_VDBB.scala 97:17:@9189.4]
  assign TPU_2_io_in_A_1_1 = 32'sh0; // @[STA_VDBB.scala 97:17:@9190.4]
  assign TPU_2_io_in_A_1_2 = 32'sh0; // @[STA_VDBB.scala 97:17:@9191.4]
  assign TPU_2_io_in_A_1_3 = 32'sh0; // @[STA_VDBB.scala 97:17:@9192.4]
  assign TPU_2_io_in_A_1_4 = 32'sh0; // @[STA_VDBB.scala 97:17:@9193.4]
  assign TPU_2_io_in_A_1_5 = 32'sh0; // @[STA_VDBB.scala 97:17:@9194.4]
  assign TPU_2_io_in_A_1_6 = 32'sh0; // @[STA_VDBB.scala 97:17:@9195.4]
  assign TPU_2_io_in_A_1_7 = 32'sh0; // @[STA_VDBB.scala 97:17:@9196.4]
  assign TPU_2_io_in_B_0_0 = _T_43000 ? $signed(TPUs_0_out_B_0_0) : $signed(_GEN_1142); // @[STA_VDBB.scala 97:17:@9149.4]
  assign TPU_2_io_in_B_0_1 = _T_43000 ? $signed(TPUs_0_out_B_0_1) : $signed(_GEN_1143); // @[STA_VDBB.scala 97:17:@9150.4]
  assign TPU_2_io_in_B_0_2 = _T_43000 ? $signed(TPUs_0_out_B_0_2) : $signed(_GEN_1144); // @[STA_VDBB.scala 97:17:@9151.4]
  assign TPU_2_io_in_B_0_3 = _T_43000 ? $signed(TPUs_0_out_B_0_3) : $signed(_GEN_1145); // @[STA_VDBB.scala 97:17:@9152.4]
  assign TPU_2_io_in_B_0_4 = _T_43000 ? $signed(TPUs_0_out_B_0_4) : $signed(_GEN_1146); // @[STA_VDBB.scala 97:17:@9153.4]
  assign TPU_2_io_in_B_0_5 = _T_43000 ? $signed(TPUs_0_out_B_0_5) : $signed(_GEN_1147); // @[STA_VDBB.scala 97:17:@9154.4]
  assign TPU_2_io_in_B_0_6 = _T_43000 ? $signed(TPUs_0_out_B_0_6) : $signed(_GEN_1148); // @[STA_VDBB.scala 97:17:@9155.4]
  assign TPU_2_io_in_B_0_7 = _T_43000 ? $signed(TPUs_0_out_B_0_7) : $signed(_GEN_1149); // @[STA_VDBB.scala 97:17:@9156.4]
  assign TPU_2_io_in_B_1_0 = _T_43000 ? $signed(TPUs_0_out_B_1_0) : $signed(_GEN_1150); // @[STA_VDBB.scala 97:17:@9157.4]
  assign TPU_2_io_in_B_1_1 = _T_43000 ? $signed(TPUs_0_out_B_1_1) : $signed(_GEN_1151); // @[STA_VDBB.scala 97:17:@9158.4]
  assign TPU_2_io_in_B_1_2 = _T_43000 ? $signed(TPUs_0_out_B_1_2) : $signed(_GEN_1152); // @[STA_VDBB.scala 97:17:@9159.4]
  assign TPU_2_io_in_B_1_3 = _T_43000 ? $signed(TPUs_0_out_B_1_3) : $signed(_GEN_1153); // @[STA_VDBB.scala 97:17:@9160.4]
  assign TPU_2_io_in_B_1_4 = _T_43000 ? $signed(TPUs_0_out_B_1_4) : $signed(_GEN_1154); // @[STA_VDBB.scala 97:17:@9161.4]
  assign TPU_2_io_in_B_1_5 = _T_43000 ? $signed(TPUs_0_out_B_1_5) : $signed(_GEN_1155); // @[STA_VDBB.scala 97:17:@9162.4]
  assign TPU_2_io_in_B_1_6 = _T_43000 ? $signed(TPUs_0_out_B_1_6) : $signed(_GEN_1156); // @[STA_VDBB.scala 97:17:@9163.4]
  assign TPU_2_io_in_B_1_7 = _T_43000 ? $signed(TPUs_0_out_B_1_7) : $signed(_GEN_1157); // @[STA_VDBB.scala 97:17:@9164.4]
  assign TPU_2_io_in_B_2_0 = _T_43000 ? $signed(TPUs_0_out_B_2_0) : $signed(_GEN_1158); // @[STA_VDBB.scala 97:17:@9165.4]
  assign TPU_2_io_in_B_2_1 = _T_43000 ? $signed(TPUs_0_out_B_2_1) : $signed(_GEN_1159); // @[STA_VDBB.scala 97:17:@9166.4]
  assign TPU_2_io_in_B_2_2 = _T_43000 ? $signed(TPUs_0_out_B_2_2) : $signed(_GEN_1160); // @[STA_VDBB.scala 97:17:@9167.4]
  assign TPU_2_io_in_B_2_3 = _T_43000 ? $signed(TPUs_0_out_B_2_3) : $signed(_GEN_1161); // @[STA_VDBB.scala 97:17:@9168.4]
  assign TPU_2_io_in_B_2_4 = _T_43000 ? $signed(TPUs_0_out_B_2_4) : $signed(_GEN_1162); // @[STA_VDBB.scala 97:17:@9169.4]
  assign TPU_2_io_in_B_2_5 = _T_43000 ? $signed(TPUs_0_out_B_2_5) : $signed(_GEN_1163); // @[STA_VDBB.scala 97:17:@9170.4]
  assign TPU_2_io_in_B_2_6 = _T_43000 ? $signed(TPUs_0_out_B_2_6) : $signed(_GEN_1164); // @[STA_VDBB.scala 97:17:@9171.4]
  assign TPU_2_io_in_B_2_7 = _T_43000 ? $signed(TPUs_0_out_B_2_7) : $signed(_GEN_1165); // @[STA_VDBB.scala 97:17:@9172.4]
  assign TPU_2_io_in_B_3_0 = _T_43000 ? $signed(TPUs_0_out_B_3_0) : $signed(_GEN_1166); // @[STA_VDBB.scala 97:17:@9173.4]
  assign TPU_2_io_in_B_3_1 = _T_43000 ? $signed(TPUs_0_out_B_3_1) : $signed(_GEN_1167); // @[STA_VDBB.scala 97:17:@9174.4]
  assign TPU_2_io_in_B_3_2 = _T_43000 ? $signed(TPUs_0_out_B_3_2) : $signed(_GEN_1168); // @[STA_VDBB.scala 97:17:@9175.4]
  assign TPU_2_io_in_B_3_3 = _T_43000 ? $signed(TPUs_0_out_B_3_3) : $signed(_GEN_1169); // @[STA_VDBB.scala 97:17:@9176.4]
  assign TPU_2_io_in_B_3_4 = _T_43000 ? $signed(TPUs_0_out_B_3_4) : $signed(_GEN_1170); // @[STA_VDBB.scala 97:17:@9177.4]
  assign TPU_2_io_in_B_3_5 = _T_43000 ? $signed(TPUs_0_out_B_3_5) : $signed(_GEN_1171); // @[STA_VDBB.scala 97:17:@9178.4]
  assign TPU_2_io_in_B_3_6 = _T_43000 ? $signed(TPUs_0_out_B_3_6) : $signed(_GEN_1172); // @[STA_VDBB.scala 97:17:@9179.4]
  assign TPU_2_io_in_B_3_7 = _T_43000 ? $signed(TPUs_0_out_B_3_7) : $signed(_GEN_1173); // @[STA_VDBB.scala 97:17:@9180.4]
  assign TPU_2_io_in_tag_0_0 = _T_43000 ? TPUs_0_out_tag_0_0 : _GEN_1174; // @[STA_VDBB.scala 97:17:@9117.4]
  assign TPU_2_io_in_tag_0_1 = _T_43000 ? TPUs_0_out_tag_0_1 : _GEN_1175; // @[STA_VDBB.scala 97:17:@9118.4]
  assign TPU_2_io_in_tag_0_2 = _T_43000 ? TPUs_0_out_tag_0_2 : _GEN_1176; // @[STA_VDBB.scala 97:17:@9119.4]
  assign TPU_2_io_in_tag_0_3 = _T_43000 ? TPUs_0_out_tag_0_3 : _GEN_1177; // @[STA_VDBB.scala 97:17:@9120.4]
  assign TPU_2_io_in_tag_0_4 = _T_43000 ? TPUs_0_out_tag_0_4 : _GEN_1178; // @[STA_VDBB.scala 97:17:@9121.4]
  assign TPU_2_io_in_tag_0_5 = _T_43000 ? TPUs_0_out_tag_0_5 : _GEN_1179; // @[STA_VDBB.scala 97:17:@9122.4]
  assign TPU_2_io_in_tag_0_6 = _T_43000 ? TPUs_0_out_tag_0_6 : _GEN_1180; // @[STA_VDBB.scala 97:17:@9123.4]
  assign TPU_2_io_in_tag_0_7 = _T_43000 ? TPUs_0_out_tag_0_7 : _GEN_1181; // @[STA_VDBB.scala 97:17:@9124.4]
  assign TPU_2_io_in_tag_1_0 = _T_43000 ? TPUs_0_out_tag_1_0 : _GEN_1182; // @[STA_VDBB.scala 97:17:@9125.4]
  assign TPU_2_io_in_tag_1_1 = _T_43000 ? TPUs_0_out_tag_1_1 : _GEN_1183; // @[STA_VDBB.scala 97:17:@9126.4]
  assign TPU_2_io_in_tag_1_2 = _T_43000 ? TPUs_0_out_tag_1_2 : _GEN_1184; // @[STA_VDBB.scala 97:17:@9127.4]
  assign TPU_2_io_in_tag_1_3 = _T_43000 ? TPUs_0_out_tag_1_3 : _GEN_1185; // @[STA_VDBB.scala 97:17:@9128.4]
  assign TPU_2_io_in_tag_1_4 = _T_43000 ? TPUs_0_out_tag_1_4 : _GEN_1186; // @[STA_VDBB.scala 97:17:@9129.4]
  assign TPU_2_io_in_tag_1_5 = _T_43000 ? TPUs_0_out_tag_1_5 : _GEN_1187; // @[STA_VDBB.scala 97:17:@9130.4]
  assign TPU_2_io_in_tag_1_6 = _T_43000 ? TPUs_0_out_tag_1_6 : _GEN_1188; // @[STA_VDBB.scala 97:17:@9131.4]
  assign TPU_2_io_in_tag_1_7 = _T_43000 ? TPUs_0_out_tag_1_7 : _GEN_1189; // @[STA_VDBB.scala 97:17:@9132.4]
  assign TPU_2_io_in_tag_2_0 = _T_43000 ? TPUs_0_out_tag_2_0 : _GEN_1190; // @[STA_VDBB.scala 97:17:@9133.4]
  assign TPU_2_io_in_tag_2_1 = _T_43000 ? TPUs_0_out_tag_2_1 : _GEN_1191; // @[STA_VDBB.scala 97:17:@9134.4]
  assign TPU_2_io_in_tag_2_2 = _T_43000 ? TPUs_0_out_tag_2_2 : _GEN_1192; // @[STA_VDBB.scala 97:17:@9135.4]
  assign TPU_2_io_in_tag_2_3 = _T_43000 ? TPUs_0_out_tag_2_3 : _GEN_1193; // @[STA_VDBB.scala 97:17:@9136.4]
  assign TPU_2_io_in_tag_2_4 = _T_43000 ? TPUs_0_out_tag_2_4 : _GEN_1194; // @[STA_VDBB.scala 97:17:@9137.4]
  assign TPU_2_io_in_tag_2_5 = _T_43000 ? TPUs_0_out_tag_2_5 : _GEN_1195; // @[STA_VDBB.scala 97:17:@9138.4]
  assign TPU_2_io_in_tag_2_6 = _T_43000 ? TPUs_0_out_tag_2_6 : _GEN_1196; // @[STA_VDBB.scala 97:17:@9139.4]
  assign TPU_2_io_in_tag_2_7 = _T_43000 ? TPUs_0_out_tag_2_7 : _GEN_1197; // @[STA_VDBB.scala 97:17:@9140.4]
  assign TPU_2_io_in_tag_3_0 = _T_43000 ? TPUs_0_out_tag_3_0 : _GEN_1198; // @[STA_VDBB.scala 97:17:@9141.4]
  assign TPU_2_io_in_tag_3_1 = _T_43000 ? TPUs_0_out_tag_3_1 : _GEN_1199; // @[STA_VDBB.scala 97:17:@9142.4]
  assign TPU_2_io_in_tag_3_2 = _T_43000 ? TPUs_0_out_tag_3_2 : _GEN_1200; // @[STA_VDBB.scala 97:17:@9143.4]
  assign TPU_2_io_in_tag_3_3 = _T_43000 ? TPUs_0_out_tag_3_3 : _GEN_1201; // @[STA_VDBB.scala 97:17:@9144.4]
  assign TPU_2_io_in_tag_3_4 = _T_43000 ? TPUs_0_out_tag_3_4 : _GEN_1202; // @[STA_VDBB.scala 97:17:@9145.4]
  assign TPU_2_io_in_tag_3_5 = _T_43000 ? TPUs_0_out_tag_3_5 : _GEN_1203; // @[STA_VDBB.scala 97:17:@9146.4]
  assign TPU_2_io_in_tag_3_6 = _T_43000 ? TPUs_0_out_tag_3_6 : _GEN_1204; // @[STA_VDBB.scala 97:17:@9147.4]
  assign TPU_2_io_in_tag_3_7 = _T_43000 ? TPUs_0_out_tag_3_7 : _GEN_1205; // @[STA_VDBB.scala 97:17:@9148.4]
  assign TPU_2_io_in_cal = cal_control_1; // @[STA_VDBB.scala 97:17:@9116.4]
  assign TPU_3_clock = clock; // @[:@8684.4]
  assign TPU_3_reset = reset; // @[:@8685.4]
  assign TPU_3_io_in_A_0_0 = TPU_2_io_out_A_0_0; // @[STA_VDBB.scala 97:17:@9351.4]
  assign TPU_3_io_in_A_0_1 = TPU_2_io_out_A_0_1; // @[STA_VDBB.scala 97:17:@9352.4]
  assign TPU_3_io_in_A_0_2 = TPU_2_io_out_A_0_2; // @[STA_VDBB.scala 97:17:@9353.4]
  assign TPU_3_io_in_A_0_3 = TPU_2_io_out_A_0_3; // @[STA_VDBB.scala 97:17:@9354.4]
  assign TPU_3_io_in_A_0_4 = TPU_2_io_out_A_0_4; // @[STA_VDBB.scala 97:17:@9355.4]
  assign TPU_3_io_in_A_0_5 = TPU_2_io_out_A_0_5; // @[STA_VDBB.scala 97:17:@9356.4]
  assign TPU_3_io_in_A_0_6 = TPU_2_io_out_A_0_6; // @[STA_VDBB.scala 97:17:@9357.4]
  assign TPU_3_io_in_A_0_7 = TPU_2_io_out_A_0_7; // @[STA_VDBB.scala 97:17:@9358.4]
  assign TPU_3_io_in_A_1_0 = TPU_2_io_out_A_1_0; // @[STA_VDBB.scala 97:17:@9359.4]
  assign TPU_3_io_in_A_1_1 = TPU_2_io_out_A_1_1; // @[STA_VDBB.scala 97:17:@9360.4]
  assign TPU_3_io_in_A_1_2 = TPU_2_io_out_A_1_2; // @[STA_VDBB.scala 97:17:@9361.4]
  assign TPU_3_io_in_A_1_3 = TPU_2_io_out_A_1_3; // @[STA_VDBB.scala 97:17:@9362.4]
  assign TPU_3_io_in_A_1_4 = TPU_2_io_out_A_1_4; // @[STA_VDBB.scala 97:17:@9363.4]
  assign TPU_3_io_in_A_1_5 = TPU_2_io_out_A_1_5; // @[STA_VDBB.scala 97:17:@9364.4]
  assign TPU_3_io_in_A_1_6 = TPU_2_io_out_A_1_6; // @[STA_VDBB.scala 97:17:@9365.4]
  assign TPU_3_io_in_A_1_7 = TPU_2_io_out_A_1_7; // @[STA_VDBB.scala 97:17:@9366.4]
  assign TPU_3_io_in_B_0_0 = TPU_1_io_out_B_0_0; // @[STA_VDBB.scala 97:17:@9319.4]
  assign TPU_3_io_in_B_0_1 = TPU_1_io_out_B_0_1; // @[STA_VDBB.scala 97:17:@9320.4]
  assign TPU_3_io_in_B_0_2 = TPU_1_io_out_B_0_2; // @[STA_VDBB.scala 97:17:@9321.4]
  assign TPU_3_io_in_B_0_3 = TPU_1_io_out_B_0_3; // @[STA_VDBB.scala 97:17:@9322.4]
  assign TPU_3_io_in_B_0_4 = TPU_1_io_out_B_0_4; // @[STA_VDBB.scala 97:17:@9323.4]
  assign TPU_3_io_in_B_0_5 = TPU_1_io_out_B_0_5; // @[STA_VDBB.scala 97:17:@9324.4]
  assign TPU_3_io_in_B_0_6 = TPU_1_io_out_B_0_6; // @[STA_VDBB.scala 97:17:@9325.4]
  assign TPU_3_io_in_B_0_7 = TPU_1_io_out_B_0_7; // @[STA_VDBB.scala 97:17:@9326.4]
  assign TPU_3_io_in_B_1_0 = TPU_1_io_out_B_1_0; // @[STA_VDBB.scala 97:17:@9327.4]
  assign TPU_3_io_in_B_1_1 = TPU_1_io_out_B_1_1; // @[STA_VDBB.scala 97:17:@9328.4]
  assign TPU_3_io_in_B_1_2 = TPU_1_io_out_B_1_2; // @[STA_VDBB.scala 97:17:@9329.4]
  assign TPU_3_io_in_B_1_3 = TPU_1_io_out_B_1_3; // @[STA_VDBB.scala 97:17:@9330.4]
  assign TPU_3_io_in_B_1_4 = TPU_1_io_out_B_1_4; // @[STA_VDBB.scala 97:17:@9331.4]
  assign TPU_3_io_in_B_1_5 = TPU_1_io_out_B_1_5; // @[STA_VDBB.scala 97:17:@9332.4]
  assign TPU_3_io_in_B_1_6 = TPU_1_io_out_B_1_6; // @[STA_VDBB.scala 97:17:@9333.4]
  assign TPU_3_io_in_B_1_7 = TPU_1_io_out_B_1_7; // @[STA_VDBB.scala 97:17:@9334.4]
  assign TPU_3_io_in_B_2_0 = TPU_1_io_out_B_2_0; // @[STA_VDBB.scala 97:17:@9335.4]
  assign TPU_3_io_in_B_2_1 = TPU_1_io_out_B_2_1; // @[STA_VDBB.scala 97:17:@9336.4]
  assign TPU_3_io_in_B_2_2 = TPU_1_io_out_B_2_2; // @[STA_VDBB.scala 97:17:@9337.4]
  assign TPU_3_io_in_B_2_3 = TPU_1_io_out_B_2_3; // @[STA_VDBB.scala 97:17:@9338.4]
  assign TPU_3_io_in_B_2_4 = TPU_1_io_out_B_2_4; // @[STA_VDBB.scala 97:17:@9339.4]
  assign TPU_3_io_in_B_2_5 = TPU_1_io_out_B_2_5; // @[STA_VDBB.scala 97:17:@9340.4]
  assign TPU_3_io_in_B_2_6 = TPU_1_io_out_B_2_6; // @[STA_VDBB.scala 97:17:@9341.4]
  assign TPU_3_io_in_B_2_7 = TPU_1_io_out_B_2_7; // @[STA_VDBB.scala 97:17:@9342.4]
  assign TPU_3_io_in_B_3_0 = TPU_1_io_out_B_3_0; // @[STA_VDBB.scala 97:17:@9343.4]
  assign TPU_3_io_in_B_3_1 = TPU_1_io_out_B_3_1; // @[STA_VDBB.scala 97:17:@9344.4]
  assign TPU_3_io_in_B_3_2 = TPU_1_io_out_B_3_2; // @[STA_VDBB.scala 97:17:@9345.4]
  assign TPU_3_io_in_B_3_3 = TPU_1_io_out_B_3_3; // @[STA_VDBB.scala 97:17:@9346.4]
  assign TPU_3_io_in_B_3_4 = TPU_1_io_out_B_3_4; // @[STA_VDBB.scala 97:17:@9347.4]
  assign TPU_3_io_in_B_3_5 = TPU_1_io_out_B_3_5; // @[STA_VDBB.scala 97:17:@9348.4]
  assign TPU_3_io_in_B_3_6 = TPU_1_io_out_B_3_6; // @[STA_VDBB.scala 97:17:@9349.4]
  assign TPU_3_io_in_B_3_7 = TPU_1_io_out_B_3_7; // @[STA_VDBB.scala 97:17:@9350.4]
  assign TPU_3_io_in_tag_0_0 = TPU_1_io_out_tag_0_0; // @[STA_VDBB.scala 97:17:@9287.4]
  assign TPU_3_io_in_tag_0_1 = TPU_1_io_out_tag_0_1; // @[STA_VDBB.scala 97:17:@9288.4]
  assign TPU_3_io_in_tag_0_2 = TPU_1_io_out_tag_0_2; // @[STA_VDBB.scala 97:17:@9289.4]
  assign TPU_3_io_in_tag_0_3 = TPU_1_io_out_tag_0_3; // @[STA_VDBB.scala 97:17:@9290.4]
  assign TPU_3_io_in_tag_0_4 = TPU_1_io_out_tag_0_4; // @[STA_VDBB.scala 97:17:@9291.4]
  assign TPU_3_io_in_tag_0_5 = TPU_1_io_out_tag_0_5; // @[STA_VDBB.scala 97:17:@9292.4]
  assign TPU_3_io_in_tag_0_6 = TPU_1_io_out_tag_0_6; // @[STA_VDBB.scala 97:17:@9293.4]
  assign TPU_3_io_in_tag_0_7 = TPU_1_io_out_tag_0_7; // @[STA_VDBB.scala 97:17:@9294.4]
  assign TPU_3_io_in_tag_1_0 = TPU_1_io_out_tag_1_0; // @[STA_VDBB.scala 97:17:@9295.4]
  assign TPU_3_io_in_tag_1_1 = TPU_1_io_out_tag_1_1; // @[STA_VDBB.scala 97:17:@9296.4]
  assign TPU_3_io_in_tag_1_2 = TPU_1_io_out_tag_1_2; // @[STA_VDBB.scala 97:17:@9297.4]
  assign TPU_3_io_in_tag_1_3 = TPU_1_io_out_tag_1_3; // @[STA_VDBB.scala 97:17:@9298.4]
  assign TPU_3_io_in_tag_1_4 = TPU_1_io_out_tag_1_4; // @[STA_VDBB.scala 97:17:@9299.4]
  assign TPU_3_io_in_tag_1_5 = TPU_1_io_out_tag_1_5; // @[STA_VDBB.scala 97:17:@9300.4]
  assign TPU_3_io_in_tag_1_6 = TPU_1_io_out_tag_1_6; // @[STA_VDBB.scala 97:17:@9301.4]
  assign TPU_3_io_in_tag_1_7 = TPU_1_io_out_tag_1_7; // @[STA_VDBB.scala 97:17:@9302.4]
  assign TPU_3_io_in_tag_2_0 = TPU_1_io_out_tag_2_0; // @[STA_VDBB.scala 97:17:@9303.4]
  assign TPU_3_io_in_tag_2_1 = TPU_1_io_out_tag_2_1; // @[STA_VDBB.scala 97:17:@9304.4]
  assign TPU_3_io_in_tag_2_2 = TPU_1_io_out_tag_2_2; // @[STA_VDBB.scala 97:17:@9305.4]
  assign TPU_3_io_in_tag_2_3 = TPU_1_io_out_tag_2_3; // @[STA_VDBB.scala 97:17:@9306.4]
  assign TPU_3_io_in_tag_2_4 = TPU_1_io_out_tag_2_4; // @[STA_VDBB.scala 97:17:@9307.4]
  assign TPU_3_io_in_tag_2_5 = TPU_1_io_out_tag_2_5; // @[STA_VDBB.scala 97:17:@9308.4]
  assign TPU_3_io_in_tag_2_6 = TPU_1_io_out_tag_2_6; // @[STA_VDBB.scala 97:17:@9309.4]
  assign TPU_3_io_in_tag_2_7 = TPU_1_io_out_tag_2_7; // @[STA_VDBB.scala 97:17:@9310.4]
  assign TPU_3_io_in_tag_3_0 = TPU_1_io_out_tag_3_0; // @[STA_VDBB.scala 97:17:@9311.4]
  assign TPU_3_io_in_tag_3_1 = TPU_1_io_out_tag_3_1; // @[STA_VDBB.scala 97:17:@9312.4]
  assign TPU_3_io_in_tag_3_2 = TPU_1_io_out_tag_3_2; // @[STA_VDBB.scala 97:17:@9313.4]
  assign TPU_3_io_in_tag_3_3 = TPU_1_io_out_tag_3_3; // @[STA_VDBB.scala 97:17:@9314.4]
  assign TPU_3_io_in_tag_3_4 = TPU_1_io_out_tag_3_4; // @[STA_VDBB.scala 97:17:@9315.4]
  assign TPU_3_io_in_tag_3_5 = TPU_1_io_out_tag_3_5; // @[STA_VDBB.scala 97:17:@9316.4]
  assign TPU_3_io_in_tag_3_6 = TPU_1_io_out_tag_3_6; // @[STA_VDBB.scala 97:17:@9317.4]
  assign TPU_3_io_in_tag_3_7 = TPU_1_io_out_tag_3_7; // @[STA_VDBB.scala 97:17:@9318.4]
  assign TPU_3_io_in_cal = cal_control_2; // @[STA_VDBB.scala 97:17:@9286.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
    `ifndef verilator
      #0.002 begin end
    `endif
  `ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  reg_A_1_0_0 = _RAND_0[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  reg_A_1_0_1 = _RAND_1[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  reg_A_1_0_2 = _RAND_2[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  reg_A_1_0_3 = _RAND_3[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  reg_A_1_0_4 = _RAND_4[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  reg_A_1_0_5 = _RAND_5[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  reg_A_1_0_6 = _RAND_6[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  reg_A_1_0_7 = _RAND_7[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  reg_A_1_1_0 = _RAND_8[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  reg_A_1_1_1 = _RAND_9[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  reg_A_1_1_2 = _RAND_10[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  reg_A_1_1_3 = _RAND_11[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  reg_A_1_1_4 = _RAND_12[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  reg_A_1_1_5 = _RAND_13[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  reg_A_1_1_6 = _RAND_14[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  reg_A_1_1_7 = _RAND_15[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  reg_A_2_0_0 = _RAND_16[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  reg_A_2_0_1 = _RAND_17[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  reg_A_2_0_2 = _RAND_18[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  reg_A_2_0_3 = _RAND_19[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  reg_A_2_0_4 = _RAND_20[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  reg_A_2_0_5 = _RAND_21[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  reg_A_2_0_6 = _RAND_22[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  reg_A_2_0_7 = _RAND_23[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  reg_A_2_1_0 = _RAND_24[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  reg_A_2_1_1 = _RAND_25[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  reg_A_2_1_2 = _RAND_26[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  reg_A_2_1_3 = _RAND_27[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  reg_A_2_1_4 = _RAND_28[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  reg_A_2_1_5 = _RAND_29[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  reg_A_2_1_6 = _RAND_30[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  reg_A_2_1_7 = _RAND_31[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  reg_A_3_0_0 = _RAND_32[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  reg_A_3_0_1 = _RAND_33[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  reg_A_3_0_2 = _RAND_34[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  reg_A_3_0_3 = _RAND_35[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  reg_A_3_0_4 = _RAND_36[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  reg_A_3_0_5 = _RAND_37[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  reg_A_3_0_6 = _RAND_38[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  reg_A_3_0_7 = _RAND_39[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  reg_A_3_1_0 = _RAND_40[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  reg_A_3_1_1 = _RAND_41[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  reg_A_3_1_2 = _RAND_42[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  reg_A_3_1_3 = _RAND_43[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  reg_A_3_1_4 = _RAND_44[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  reg_A_3_1_5 = _RAND_45[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  reg_A_3_1_6 = _RAND_46[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  reg_A_3_1_7 = _RAND_47[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  reg_A_4_0_0 = _RAND_48[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  reg_A_4_0_1 = _RAND_49[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  reg_A_4_0_2 = _RAND_50[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  reg_A_4_0_3 = _RAND_51[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  reg_A_4_0_4 = _RAND_52[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  reg_A_4_0_5 = _RAND_53[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  reg_A_4_0_6 = _RAND_54[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  reg_A_4_0_7 = _RAND_55[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  reg_A_4_1_0 = _RAND_56[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  reg_A_4_1_1 = _RAND_57[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  reg_A_4_1_2 = _RAND_58[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  reg_A_4_1_3 = _RAND_59[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  reg_A_4_1_4 = _RAND_60[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  reg_A_4_1_5 = _RAND_61[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  reg_A_4_1_6 = _RAND_62[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  reg_A_4_1_7 = _RAND_63[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_64 = {1{$random}};
  reg_B_1_0_0 = _RAND_64[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_65 = {1{$random}};
  reg_B_1_0_1 = _RAND_65[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_66 = {1{$random}};
  reg_B_1_0_2 = _RAND_66[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_67 = {1{$random}};
  reg_B_1_0_3 = _RAND_67[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_68 = {1{$random}};
  reg_B_1_0_4 = _RAND_68[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_69 = {1{$random}};
  reg_B_1_0_5 = _RAND_69[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_70 = {1{$random}};
  reg_B_1_0_6 = _RAND_70[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_71 = {1{$random}};
  reg_B_1_0_7 = _RAND_71[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_72 = {1{$random}};
  reg_B_1_1_0 = _RAND_72[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_73 = {1{$random}};
  reg_B_1_1_1 = _RAND_73[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_74 = {1{$random}};
  reg_B_1_1_2 = _RAND_74[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_75 = {1{$random}};
  reg_B_1_1_3 = _RAND_75[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_76 = {1{$random}};
  reg_B_1_1_4 = _RAND_76[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_77 = {1{$random}};
  reg_B_1_1_5 = _RAND_77[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_78 = {1{$random}};
  reg_B_1_1_6 = _RAND_78[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_79 = {1{$random}};
  reg_B_1_1_7 = _RAND_79[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_80 = {1{$random}};
  reg_B_1_2_0 = _RAND_80[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_81 = {1{$random}};
  reg_B_1_2_1 = _RAND_81[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_82 = {1{$random}};
  reg_B_1_2_2 = _RAND_82[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_83 = {1{$random}};
  reg_B_1_2_3 = _RAND_83[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_84 = {1{$random}};
  reg_B_1_2_4 = _RAND_84[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_85 = {1{$random}};
  reg_B_1_2_5 = _RAND_85[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_86 = {1{$random}};
  reg_B_1_2_6 = _RAND_86[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_87 = {1{$random}};
  reg_B_1_2_7 = _RAND_87[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_88 = {1{$random}};
  reg_B_1_3_0 = _RAND_88[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_89 = {1{$random}};
  reg_B_1_3_1 = _RAND_89[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_90 = {1{$random}};
  reg_B_1_3_2 = _RAND_90[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_91 = {1{$random}};
  reg_B_1_3_3 = _RAND_91[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_92 = {1{$random}};
  reg_B_1_3_4 = _RAND_92[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_93 = {1{$random}};
  reg_B_1_3_5 = _RAND_93[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_94 = {1{$random}};
  reg_B_1_3_6 = _RAND_94[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_95 = {1{$random}};
  reg_B_1_3_7 = _RAND_95[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_96 = {1{$random}};
  reg_B_2_0_0 = _RAND_96[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_97 = {1{$random}};
  reg_B_2_0_1 = _RAND_97[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_98 = {1{$random}};
  reg_B_2_0_2 = _RAND_98[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_99 = {1{$random}};
  reg_B_2_0_3 = _RAND_99[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_100 = {1{$random}};
  reg_B_2_0_4 = _RAND_100[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_101 = {1{$random}};
  reg_B_2_0_5 = _RAND_101[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_102 = {1{$random}};
  reg_B_2_0_6 = _RAND_102[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_103 = {1{$random}};
  reg_B_2_0_7 = _RAND_103[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_104 = {1{$random}};
  reg_B_2_1_0 = _RAND_104[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_105 = {1{$random}};
  reg_B_2_1_1 = _RAND_105[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_106 = {1{$random}};
  reg_B_2_1_2 = _RAND_106[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_107 = {1{$random}};
  reg_B_2_1_3 = _RAND_107[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_108 = {1{$random}};
  reg_B_2_1_4 = _RAND_108[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_109 = {1{$random}};
  reg_B_2_1_5 = _RAND_109[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_110 = {1{$random}};
  reg_B_2_1_6 = _RAND_110[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_111 = {1{$random}};
  reg_B_2_1_7 = _RAND_111[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_112 = {1{$random}};
  reg_B_2_2_0 = _RAND_112[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_113 = {1{$random}};
  reg_B_2_2_1 = _RAND_113[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_114 = {1{$random}};
  reg_B_2_2_2 = _RAND_114[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_115 = {1{$random}};
  reg_B_2_2_3 = _RAND_115[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_116 = {1{$random}};
  reg_B_2_2_4 = _RAND_116[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_117 = {1{$random}};
  reg_B_2_2_5 = _RAND_117[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_118 = {1{$random}};
  reg_B_2_2_6 = _RAND_118[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_119 = {1{$random}};
  reg_B_2_2_7 = _RAND_119[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_120 = {1{$random}};
  reg_B_2_3_0 = _RAND_120[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_121 = {1{$random}};
  reg_B_2_3_1 = _RAND_121[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_122 = {1{$random}};
  reg_B_2_3_2 = _RAND_122[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_123 = {1{$random}};
  reg_B_2_3_3 = _RAND_123[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_124 = {1{$random}};
  reg_B_2_3_4 = _RAND_124[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_125 = {1{$random}};
  reg_B_2_3_5 = _RAND_125[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_126 = {1{$random}};
  reg_B_2_3_6 = _RAND_126[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_127 = {1{$random}};
  reg_B_2_3_7 = _RAND_127[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_128 = {1{$random}};
  reg_B_3_0_0 = _RAND_128[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_129 = {1{$random}};
  reg_B_3_0_1 = _RAND_129[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_130 = {1{$random}};
  reg_B_3_0_2 = _RAND_130[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_131 = {1{$random}};
  reg_B_3_0_3 = _RAND_131[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_132 = {1{$random}};
  reg_B_3_0_4 = _RAND_132[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_133 = {1{$random}};
  reg_B_3_0_5 = _RAND_133[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_134 = {1{$random}};
  reg_B_3_0_6 = _RAND_134[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_135 = {1{$random}};
  reg_B_3_0_7 = _RAND_135[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_136 = {1{$random}};
  reg_B_3_1_0 = _RAND_136[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_137 = {1{$random}};
  reg_B_3_1_1 = _RAND_137[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_138 = {1{$random}};
  reg_B_3_1_2 = _RAND_138[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_139 = {1{$random}};
  reg_B_3_1_3 = _RAND_139[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_140 = {1{$random}};
  reg_B_3_1_4 = _RAND_140[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_141 = {1{$random}};
  reg_B_3_1_5 = _RAND_141[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_142 = {1{$random}};
  reg_B_3_1_6 = _RAND_142[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_143 = {1{$random}};
  reg_B_3_1_7 = _RAND_143[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_144 = {1{$random}};
  reg_B_3_2_0 = _RAND_144[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_145 = {1{$random}};
  reg_B_3_2_1 = _RAND_145[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_146 = {1{$random}};
  reg_B_3_2_2 = _RAND_146[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_147 = {1{$random}};
  reg_B_3_2_3 = _RAND_147[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_148 = {1{$random}};
  reg_B_3_2_4 = _RAND_148[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_149 = {1{$random}};
  reg_B_3_2_5 = _RAND_149[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_150 = {1{$random}};
  reg_B_3_2_6 = _RAND_150[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_151 = {1{$random}};
  reg_B_3_2_7 = _RAND_151[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_152 = {1{$random}};
  reg_B_3_3_0 = _RAND_152[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_153 = {1{$random}};
  reg_B_3_3_1 = _RAND_153[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_154 = {1{$random}};
  reg_B_3_3_2 = _RAND_154[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_155 = {1{$random}};
  reg_B_3_3_3 = _RAND_155[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_156 = {1{$random}};
  reg_B_3_3_4 = _RAND_156[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_157 = {1{$random}};
  reg_B_3_3_5 = _RAND_157[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_158 = {1{$random}};
  reg_B_3_3_6 = _RAND_158[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_159 = {1{$random}};
  reg_B_3_3_7 = _RAND_159[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_160 = {1{$random}};
  reg_B_4_0_0 = _RAND_160[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_161 = {1{$random}};
  reg_B_4_0_1 = _RAND_161[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_162 = {1{$random}};
  reg_B_4_0_2 = _RAND_162[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_163 = {1{$random}};
  reg_B_4_0_3 = _RAND_163[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_164 = {1{$random}};
  reg_B_4_0_4 = _RAND_164[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_165 = {1{$random}};
  reg_B_4_0_5 = _RAND_165[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_166 = {1{$random}};
  reg_B_4_0_6 = _RAND_166[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_167 = {1{$random}};
  reg_B_4_0_7 = _RAND_167[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_168 = {1{$random}};
  reg_B_4_1_0 = _RAND_168[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_169 = {1{$random}};
  reg_B_4_1_1 = _RAND_169[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_170 = {1{$random}};
  reg_B_4_1_2 = _RAND_170[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_171 = {1{$random}};
  reg_B_4_1_3 = _RAND_171[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_172 = {1{$random}};
  reg_B_4_1_4 = _RAND_172[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_173 = {1{$random}};
  reg_B_4_1_5 = _RAND_173[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_174 = {1{$random}};
  reg_B_4_1_6 = _RAND_174[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_175 = {1{$random}};
  reg_B_4_1_7 = _RAND_175[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_176 = {1{$random}};
  reg_B_4_2_0 = _RAND_176[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_177 = {1{$random}};
  reg_B_4_2_1 = _RAND_177[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_178 = {1{$random}};
  reg_B_4_2_2 = _RAND_178[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_179 = {1{$random}};
  reg_B_4_2_3 = _RAND_179[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_180 = {1{$random}};
  reg_B_4_2_4 = _RAND_180[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_181 = {1{$random}};
  reg_B_4_2_5 = _RAND_181[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_182 = {1{$random}};
  reg_B_4_2_6 = _RAND_182[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_183 = {1{$random}};
  reg_B_4_2_7 = _RAND_183[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_184 = {1{$random}};
  reg_B_4_3_0 = _RAND_184[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_185 = {1{$random}};
  reg_B_4_3_1 = _RAND_185[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_186 = {1{$random}};
  reg_B_4_3_2 = _RAND_186[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_187 = {1{$random}};
  reg_B_4_3_3 = _RAND_187[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_188 = {1{$random}};
  reg_B_4_3_4 = _RAND_188[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_189 = {1{$random}};
  reg_B_4_3_5 = _RAND_189[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_190 = {1{$random}};
  reg_B_4_3_6 = _RAND_190[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_191 = {1{$random}};
  reg_B_4_3_7 = _RAND_191[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_192 = {1{$random}};
  cal_state_0 = _RAND_192[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_193 = {1{$random}};
  cal_state_1 = _RAND_193[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_194 = {1{$random}};
  cal_state_2 = _RAND_194[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_195 = {1{$random}};
  result_0_0 = _RAND_195[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_196 = {1{$random}};
  result_0_1 = _RAND_196[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_197 = {1{$random}};
  result_0_2 = _RAND_197[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_198 = {1{$random}};
  result_0_3 = _RAND_198[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_199 = {1{$random}};
  result_0_4 = _RAND_199[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_200 = {1{$random}};
  result_0_5 = _RAND_200[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_201 = {1{$random}};
  result_0_6 = _RAND_201[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_202 = {1{$random}};
  result_0_7 = _RAND_202[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_203 = {1{$random}};
  result_1_0 = _RAND_203[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_204 = {1{$random}};
  result_1_1 = _RAND_204[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_205 = {1{$random}};
  result_1_2 = _RAND_205[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_206 = {1{$random}};
  result_1_3 = _RAND_206[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_207 = {1{$random}};
  result_1_4 = _RAND_207[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_208 = {1{$random}};
  result_1_5 = _RAND_208[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_209 = {1{$random}};
  result_1_6 = _RAND_209[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_210 = {1{$random}};
  result_1_7 = _RAND_210[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_211 = {1{$random}};
  result_2_0 = _RAND_211[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_212 = {1{$random}};
  result_2_1 = _RAND_212[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_213 = {1{$random}};
  result_2_2 = _RAND_213[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_214 = {1{$random}};
  result_2_3 = _RAND_214[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_215 = {1{$random}};
  result_2_4 = _RAND_215[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_216 = {1{$random}};
  result_2_5 = _RAND_216[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_217 = {1{$random}};
  result_2_6 = _RAND_217[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_218 = {1{$random}};
  result_2_7 = _RAND_218[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_219 = {1{$random}};
  result_3_0 = _RAND_219[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_220 = {1{$random}};
  result_3_1 = _RAND_220[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_221 = {1{$random}};
  result_3_2 = _RAND_221[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_222 = {1{$random}};
  result_3_3 = _RAND_222[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_223 = {1{$random}};
  result_3_4 = _RAND_223[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_224 = {1{$random}};
  result_3_5 = _RAND_224[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_225 = {1{$random}};
  result_3_6 = _RAND_225[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_226 = {1{$random}};
  result_3_7 = _RAND_226[31:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_227 = {1{$random}};
  cal_control_0 = _RAND_227[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_228 = {1{$random}};
  cal_control_1 = _RAND_228[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_229 = {1{$random}};
  cal_control_2 = _RAND_229[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_230 = {1{$random}};
  stateReg = _RAND_230[2:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_231 = {1{$random}};
  loop_reg = _RAND_231[0:0];
  `endif // RANDOMIZE_REG_INIT
  `ifdef RANDOMIZE_REG_INIT
  _RAND_232 = {1{$random}};
  _T_43002 = _RAND_232[0:0];
  `endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      reg_A_1_0_0 <= 32'sh0;
    end else begin
      reg_A_1_0_0 <= io_in_A_0_0;
    end
    if (reset) begin
      reg_A_1_0_1 <= 32'sh0;
    end else begin
      reg_A_1_0_1 <= io_in_A_0_1;
    end
    if (reset) begin
      reg_A_1_0_2 <= 32'sh0;
    end else begin
      reg_A_1_0_2 <= io_in_A_0_2;
    end
    if (reset) begin
      reg_A_1_0_3 <= 32'sh0;
    end else begin
      reg_A_1_0_3 <= io_in_A_0_3;
    end
    if (reset) begin
      reg_A_1_0_4 <= 32'sh0;
    end else begin
      reg_A_1_0_4 <= io_in_A_0_4;
    end
    if (reset) begin
      reg_A_1_0_5 <= 32'sh0;
    end else begin
      reg_A_1_0_5 <= io_in_A_0_5;
    end
    if (reset) begin
      reg_A_1_0_6 <= 32'sh0;
    end else begin
      reg_A_1_0_6 <= io_in_A_0_6;
    end
    if (reset) begin
      reg_A_1_0_7 <= 32'sh0;
    end else begin
      reg_A_1_0_7 <= io_in_A_0_7;
    end
    if (reset) begin
      reg_A_1_1_0 <= 32'sh0;
    end else begin
      reg_A_1_1_0 <= io_in_A_1_0;
    end
    if (reset) begin
      reg_A_1_1_1 <= 32'sh0;
    end else begin
      reg_A_1_1_1 <= io_in_A_1_1;
    end
    if (reset) begin
      reg_A_1_1_2 <= 32'sh0;
    end else begin
      reg_A_1_1_2 <= io_in_A_1_2;
    end
    if (reset) begin
      reg_A_1_1_3 <= 32'sh0;
    end else begin
      reg_A_1_1_3 <= io_in_A_1_3;
    end
    if (reset) begin
      reg_A_1_1_4 <= 32'sh0;
    end else begin
      reg_A_1_1_4 <= io_in_A_1_4;
    end
    if (reset) begin
      reg_A_1_1_5 <= 32'sh0;
    end else begin
      reg_A_1_1_5 <= io_in_A_1_5;
    end
    if (reset) begin
      reg_A_1_1_6 <= 32'sh0;
    end else begin
      reg_A_1_1_6 <= io_in_A_1_6;
    end
    if (reset) begin
      reg_A_1_1_7 <= 32'sh0;
    end else begin
      reg_A_1_1_7 <= io_in_A_1_7;
    end
    if (reset) begin
      reg_A_2_0_0 <= 32'sh0;
    end else begin
      reg_A_2_0_0 <= io_in_A_0_8;
    end
    if (reset) begin
      reg_A_2_0_1 <= 32'sh0;
    end else begin
      reg_A_2_0_1 <= io_in_A_0_9;
    end
    if (reset) begin
      reg_A_2_0_2 <= 32'sh0;
    end else begin
      reg_A_2_0_2 <= io_in_A_0_10;
    end
    if (reset) begin
      reg_A_2_0_3 <= 32'sh0;
    end else begin
      reg_A_2_0_3 <= io_in_A_0_11;
    end
    if (reset) begin
      reg_A_2_0_4 <= 32'sh0;
    end else begin
      reg_A_2_0_4 <= io_in_A_0_12;
    end
    if (reset) begin
      reg_A_2_0_5 <= 32'sh0;
    end else begin
      reg_A_2_0_5 <= io_in_A_0_13;
    end
    if (reset) begin
      reg_A_2_0_6 <= 32'sh0;
    end else begin
      reg_A_2_0_6 <= io_in_A_0_14;
    end
    if (reset) begin
      reg_A_2_0_7 <= 32'sh0;
    end else begin
      reg_A_2_0_7 <= io_in_A_0_15;
    end
    if (reset) begin
      reg_A_2_1_0 <= 32'sh0;
    end else begin
      reg_A_2_1_0 <= io_in_A_1_8;
    end
    if (reset) begin
      reg_A_2_1_1 <= 32'sh0;
    end else begin
      reg_A_2_1_1 <= io_in_A_1_9;
    end
    if (reset) begin
      reg_A_2_1_2 <= 32'sh0;
    end else begin
      reg_A_2_1_2 <= io_in_A_1_10;
    end
    if (reset) begin
      reg_A_2_1_3 <= 32'sh0;
    end else begin
      reg_A_2_1_3 <= io_in_A_1_11;
    end
    if (reset) begin
      reg_A_2_1_4 <= 32'sh0;
    end else begin
      reg_A_2_1_4 <= io_in_A_1_12;
    end
    if (reset) begin
      reg_A_2_1_5 <= 32'sh0;
    end else begin
      reg_A_2_1_5 <= io_in_A_1_13;
    end
    if (reset) begin
      reg_A_2_1_6 <= 32'sh0;
    end else begin
      reg_A_2_1_6 <= io_in_A_1_14;
    end
    if (reset) begin
      reg_A_2_1_7 <= 32'sh0;
    end else begin
      reg_A_2_1_7 <= io_in_A_1_15;
    end
    if (reset) begin
      reg_A_3_0_0 <= 32'sh0;
    end else begin
      reg_A_3_0_0 <= io_in_A_2_0;
    end
    if (reset) begin
      reg_A_3_0_1 <= 32'sh0;
    end else begin
      reg_A_3_0_1 <= io_in_A_2_1;
    end
    if (reset) begin
      reg_A_3_0_2 <= 32'sh0;
    end else begin
      reg_A_3_0_2 <= io_in_A_2_2;
    end
    if (reset) begin
      reg_A_3_0_3 <= 32'sh0;
    end else begin
      reg_A_3_0_3 <= io_in_A_2_3;
    end
    if (reset) begin
      reg_A_3_0_4 <= 32'sh0;
    end else begin
      reg_A_3_0_4 <= io_in_A_2_4;
    end
    if (reset) begin
      reg_A_3_0_5 <= 32'sh0;
    end else begin
      reg_A_3_0_5 <= io_in_A_2_5;
    end
    if (reset) begin
      reg_A_3_0_6 <= 32'sh0;
    end else begin
      reg_A_3_0_6 <= io_in_A_2_6;
    end
    if (reset) begin
      reg_A_3_0_7 <= 32'sh0;
    end else begin
      reg_A_3_0_7 <= io_in_A_2_7;
    end
    if (reset) begin
      reg_A_3_1_0 <= 32'sh0;
    end else begin
      reg_A_3_1_0 <= io_in_A_3_0;
    end
    if (reset) begin
      reg_A_3_1_1 <= 32'sh0;
    end else begin
      reg_A_3_1_1 <= io_in_A_3_1;
    end
    if (reset) begin
      reg_A_3_1_2 <= 32'sh0;
    end else begin
      reg_A_3_1_2 <= io_in_A_3_2;
    end
    if (reset) begin
      reg_A_3_1_3 <= 32'sh0;
    end else begin
      reg_A_3_1_3 <= io_in_A_3_3;
    end
    if (reset) begin
      reg_A_3_1_4 <= 32'sh0;
    end else begin
      reg_A_3_1_4 <= io_in_A_3_4;
    end
    if (reset) begin
      reg_A_3_1_5 <= 32'sh0;
    end else begin
      reg_A_3_1_5 <= io_in_A_3_5;
    end
    if (reset) begin
      reg_A_3_1_6 <= 32'sh0;
    end else begin
      reg_A_3_1_6 <= io_in_A_3_6;
    end
    if (reset) begin
      reg_A_3_1_7 <= 32'sh0;
    end else begin
      reg_A_3_1_7 <= io_in_A_3_7;
    end
    if (reset) begin
      reg_A_4_0_0 <= 32'sh0;
    end else begin
      reg_A_4_0_0 <= io_in_A_2_8;
    end
    if (reset) begin
      reg_A_4_0_1 <= 32'sh0;
    end else begin
      reg_A_4_0_1 <= io_in_A_2_9;
    end
    if (reset) begin
      reg_A_4_0_2 <= 32'sh0;
    end else begin
      reg_A_4_0_2 <= io_in_A_2_10;
    end
    if (reset) begin
      reg_A_4_0_3 <= 32'sh0;
    end else begin
      reg_A_4_0_3 <= io_in_A_2_11;
    end
    if (reset) begin
      reg_A_4_0_4 <= 32'sh0;
    end else begin
      reg_A_4_0_4 <= io_in_A_2_12;
    end
    if (reset) begin
      reg_A_4_0_5 <= 32'sh0;
    end else begin
      reg_A_4_0_5 <= io_in_A_2_13;
    end
    if (reset) begin
      reg_A_4_0_6 <= 32'sh0;
    end else begin
      reg_A_4_0_6 <= io_in_A_2_14;
    end
    if (reset) begin
      reg_A_4_0_7 <= 32'sh0;
    end else begin
      reg_A_4_0_7 <= io_in_A_2_15;
    end
    if (reset) begin
      reg_A_4_1_0 <= 32'sh0;
    end else begin
      reg_A_4_1_0 <= io_in_A_3_8;
    end
    if (reset) begin
      reg_A_4_1_1 <= 32'sh0;
    end else begin
      reg_A_4_1_1 <= io_in_A_3_9;
    end
    if (reset) begin
      reg_A_4_1_2 <= 32'sh0;
    end else begin
      reg_A_4_1_2 <= io_in_A_3_10;
    end
    if (reset) begin
      reg_A_4_1_3 <= 32'sh0;
    end else begin
      reg_A_4_1_3 <= io_in_A_3_11;
    end
    if (reset) begin
      reg_A_4_1_4 <= 32'sh0;
    end else begin
      reg_A_4_1_4 <= io_in_A_3_12;
    end
    if (reset) begin
      reg_A_4_1_5 <= 32'sh0;
    end else begin
      reg_A_4_1_5 <= io_in_A_3_13;
    end
    if (reset) begin
      reg_A_4_1_6 <= 32'sh0;
    end else begin
      reg_A_4_1_6 <= io_in_A_3_14;
    end
    if (reset) begin
      reg_A_4_1_7 <= 32'sh0;
    end else begin
      reg_A_4_1_7 <= io_in_A_3_15;
    end
    if (reset) begin
      reg_B_1_0_0 <= 32'sh0;
    end else begin
      reg_B_1_0_0 <= io_in_B_0_0;
    end
    if (reset) begin
      reg_B_1_0_1 <= 32'sh0;
    end else begin
      reg_B_1_0_1 <= io_in_B_0_1;
    end
    if (reset) begin
      reg_B_1_0_2 <= 32'sh0;
    end else begin
      reg_B_1_0_2 <= io_in_B_0_2;
    end
    if (reset) begin
      reg_B_1_0_3 <= 32'sh0;
    end else begin
      reg_B_1_0_3 <= io_in_B_0_3;
    end
    if (reset) begin
      reg_B_1_0_4 <= 32'sh0;
    end else begin
      reg_B_1_0_4 <= io_in_B_0_4;
    end
    if (reset) begin
      reg_B_1_0_5 <= 32'sh0;
    end else begin
      reg_B_1_0_5 <= io_in_B_0_5;
    end
    if (reset) begin
      reg_B_1_0_6 <= 32'sh0;
    end else begin
      reg_B_1_0_6 <= io_in_B_0_6;
    end
    if (reset) begin
      reg_B_1_0_7 <= 32'sh0;
    end else begin
      reg_B_1_0_7 <= io_in_B_0_7;
    end
    if (reset) begin
      reg_B_1_1_0 <= 32'sh0;
    end else begin
      reg_B_1_1_0 <= io_in_B_1_0;
    end
    if (reset) begin
      reg_B_1_1_1 <= 32'sh0;
    end else begin
      reg_B_1_1_1 <= io_in_B_1_1;
    end
    if (reset) begin
      reg_B_1_1_2 <= 32'sh0;
    end else begin
      reg_B_1_1_2 <= io_in_B_1_2;
    end
    if (reset) begin
      reg_B_1_1_3 <= 32'sh0;
    end else begin
      reg_B_1_1_3 <= io_in_B_1_3;
    end
    if (reset) begin
      reg_B_1_1_4 <= 32'sh0;
    end else begin
      reg_B_1_1_4 <= io_in_B_1_4;
    end
    if (reset) begin
      reg_B_1_1_5 <= 32'sh0;
    end else begin
      reg_B_1_1_5 <= io_in_B_1_5;
    end
    if (reset) begin
      reg_B_1_1_6 <= 32'sh0;
    end else begin
      reg_B_1_1_6 <= io_in_B_1_6;
    end
    if (reset) begin
      reg_B_1_1_7 <= 32'sh0;
    end else begin
      reg_B_1_1_7 <= io_in_B_1_7;
    end
    if (reset) begin
      reg_B_1_2_0 <= 32'sh0;
    end else begin
      reg_B_1_2_0 <= io_in_B_2_0;
    end
    if (reset) begin
      reg_B_1_2_1 <= 32'sh0;
    end else begin
      reg_B_1_2_1 <= io_in_B_2_1;
    end
    if (reset) begin
      reg_B_1_2_2 <= 32'sh0;
    end else begin
      reg_B_1_2_2 <= io_in_B_2_2;
    end
    if (reset) begin
      reg_B_1_2_3 <= 32'sh0;
    end else begin
      reg_B_1_2_3 <= io_in_B_2_3;
    end
    if (reset) begin
      reg_B_1_2_4 <= 32'sh0;
    end else begin
      reg_B_1_2_4 <= io_in_B_2_4;
    end
    if (reset) begin
      reg_B_1_2_5 <= 32'sh0;
    end else begin
      reg_B_1_2_5 <= io_in_B_2_5;
    end
    if (reset) begin
      reg_B_1_2_6 <= 32'sh0;
    end else begin
      reg_B_1_2_6 <= io_in_B_2_6;
    end
    if (reset) begin
      reg_B_1_2_7 <= 32'sh0;
    end else begin
      reg_B_1_2_7 <= io_in_B_2_7;
    end
    if (reset) begin
      reg_B_1_3_0 <= 32'sh0;
    end else begin
      reg_B_1_3_0 <= io_in_B_3_0;
    end
    if (reset) begin
      reg_B_1_3_1 <= 32'sh0;
    end else begin
      reg_B_1_3_1 <= io_in_B_3_1;
    end
    if (reset) begin
      reg_B_1_3_2 <= 32'sh0;
    end else begin
      reg_B_1_3_2 <= io_in_B_3_2;
    end
    if (reset) begin
      reg_B_1_3_3 <= 32'sh0;
    end else begin
      reg_B_1_3_3 <= io_in_B_3_3;
    end
    if (reset) begin
      reg_B_1_3_4 <= 32'sh0;
    end else begin
      reg_B_1_3_4 <= io_in_B_3_4;
    end
    if (reset) begin
      reg_B_1_3_5 <= 32'sh0;
    end else begin
      reg_B_1_3_5 <= io_in_B_3_5;
    end
    if (reset) begin
      reg_B_1_3_6 <= 32'sh0;
    end else begin
      reg_B_1_3_6 <= io_in_B_3_6;
    end
    if (reset) begin
      reg_B_1_3_7 <= 32'sh0;
    end else begin
      reg_B_1_3_7 <= io_in_B_3_7;
    end
    if (reset) begin
      reg_B_2_0_0 <= 32'sh0;
    end else begin
      reg_B_2_0_0 <= io_in_B_0_8;
    end
    if (reset) begin
      reg_B_2_0_1 <= 32'sh0;
    end else begin
      reg_B_2_0_1 <= io_in_B_0_9;
    end
    if (reset) begin
      reg_B_2_0_2 <= 32'sh0;
    end else begin
      reg_B_2_0_2 <= io_in_B_0_10;
    end
    if (reset) begin
      reg_B_2_0_3 <= 32'sh0;
    end else begin
      reg_B_2_0_3 <= io_in_B_0_11;
    end
    if (reset) begin
      reg_B_2_0_4 <= 32'sh0;
    end else begin
      reg_B_2_0_4 <= io_in_B_0_12;
    end
    if (reset) begin
      reg_B_2_0_5 <= 32'sh0;
    end else begin
      reg_B_2_0_5 <= io_in_B_0_13;
    end
    if (reset) begin
      reg_B_2_0_6 <= 32'sh0;
    end else begin
      reg_B_2_0_6 <= io_in_B_0_14;
    end
    if (reset) begin
      reg_B_2_0_7 <= 32'sh0;
    end else begin
      reg_B_2_0_7 <= io_in_B_0_15;
    end
    if (reset) begin
      reg_B_2_1_0 <= 32'sh0;
    end else begin
      reg_B_2_1_0 <= io_in_B_1_8;
    end
    if (reset) begin
      reg_B_2_1_1 <= 32'sh0;
    end else begin
      reg_B_2_1_1 <= io_in_B_1_9;
    end
    if (reset) begin
      reg_B_2_1_2 <= 32'sh0;
    end else begin
      reg_B_2_1_2 <= io_in_B_1_10;
    end
    if (reset) begin
      reg_B_2_1_3 <= 32'sh0;
    end else begin
      reg_B_2_1_3 <= io_in_B_1_11;
    end
    if (reset) begin
      reg_B_2_1_4 <= 32'sh0;
    end else begin
      reg_B_2_1_4 <= io_in_B_1_12;
    end
    if (reset) begin
      reg_B_2_1_5 <= 32'sh0;
    end else begin
      reg_B_2_1_5 <= io_in_B_1_13;
    end
    if (reset) begin
      reg_B_2_1_6 <= 32'sh0;
    end else begin
      reg_B_2_1_6 <= io_in_B_1_14;
    end
    if (reset) begin
      reg_B_2_1_7 <= 32'sh0;
    end else begin
      reg_B_2_1_7 <= io_in_B_1_15;
    end
    if (reset) begin
      reg_B_2_2_0 <= 32'sh0;
    end else begin
      reg_B_2_2_0 <= io_in_B_2_8;
    end
    if (reset) begin
      reg_B_2_2_1 <= 32'sh0;
    end else begin
      reg_B_2_2_1 <= io_in_B_2_9;
    end
    if (reset) begin
      reg_B_2_2_2 <= 32'sh0;
    end else begin
      reg_B_2_2_2 <= io_in_B_2_10;
    end
    if (reset) begin
      reg_B_2_2_3 <= 32'sh0;
    end else begin
      reg_B_2_2_3 <= io_in_B_2_11;
    end
    if (reset) begin
      reg_B_2_2_4 <= 32'sh0;
    end else begin
      reg_B_2_2_4 <= io_in_B_2_12;
    end
    if (reset) begin
      reg_B_2_2_5 <= 32'sh0;
    end else begin
      reg_B_2_2_5 <= io_in_B_2_13;
    end
    if (reset) begin
      reg_B_2_2_6 <= 32'sh0;
    end else begin
      reg_B_2_2_6 <= io_in_B_2_14;
    end
    if (reset) begin
      reg_B_2_2_7 <= 32'sh0;
    end else begin
      reg_B_2_2_7 <= io_in_B_2_15;
    end
    if (reset) begin
      reg_B_2_3_0 <= 32'sh0;
    end else begin
      reg_B_2_3_0 <= io_in_B_3_8;
    end
    if (reset) begin
      reg_B_2_3_1 <= 32'sh0;
    end else begin
      reg_B_2_3_1 <= io_in_B_3_9;
    end
    if (reset) begin
      reg_B_2_3_2 <= 32'sh0;
    end else begin
      reg_B_2_3_2 <= io_in_B_3_10;
    end
    if (reset) begin
      reg_B_2_3_3 <= 32'sh0;
    end else begin
      reg_B_2_3_3 <= io_in_B_3_11;
    end
    if (reset) begin
      reg_B_2_3_4 <= 32'sh0;
    end else begin
      reg_B_2_3_4 <= io_in_B_3_12;
    end
    if (reset) begin
      reg_B_2_3_5 <= 32'sh0;
    end else begin
      reg_B_2_3_5 <= io_in_B_3_13;
    end
    if (reset) begin
      reg_B_2_3_6 <= 32'sh0;
    end else begin
      reg_B_2_3_6 <= io_in_B_3_14;
    end
    if (reset) begin
      reg_B_2_3_7 <= 32'sh0;
    end else begin
      reg_B_2_3_7 <= io_in_B_3_15;
    end
    if (reset) begin
      reg_B_3_0_0 <= 32'sh0;
    end else begin
      reg_B_3_0_0 <= io_in_B_4_0;
    end
    if (reset) begin
      reg_B_3_0_1 <= 32'sh0;
    end else begin
      reg_B_3_0_1 <= io_in_B_4_1;
    end
    if (reset) begin
      reg_B_3_0_2 <= 32'sh0;
    end else begin
      reg_B_3_0_2 <= io_in_B_4_2;
    end
    if (reset) begin
      reg_B_3_0_3 <= 32'sh0;
    end else begin
      reg_B_3_0_3 <= io_in_B_4_3;
    end
    if (reset) begin
      reg_B_3_0_4 <= 32'sh0;
    end else begin
      reg_B_3_0_4 <= io_in_B_4_4;
    end
    if (reset) begin
      reg_B_3_0_5 <= 32'sh0;
    end else begin
      reg_B_3_0_5 <= io_in_B_4_5;
    end
    if (reset) begin
      reg_B_3_0_6 <= 32'sh0;
    end else begin
      reg_B_3_0_6 <= io_in_B_4_6;
    end
    if (reset) begin
      reg_B_3_0_7 <= 32'sh0;
    end else begin
      reg_B_3_0_7 <= io_in_B_4_7;
    end
    if (reset) begin
      reg_B_3_1_0 <= 32'sh0;
    end else begin
      reg_B_3_1_0 <= io_in_B_5_0;
    end
    if (reset) begin
      reg_B_3_1_1 <= 32'sh0;
    end else begin
      reg_B_3_1_1 <= io_in_B_5_1;
    end
    if (reset) begin
      reg_B_3_1_2 <= 32'sh0;
    end else begin
      reg_B_3_1_2 <= io_in_B_5_2;
    end
    if (reset) begin
      reg_B_3_1_3 <= 32'sh0;
    end else begin
      reg_B_3_1_3 <= io_in_B_5_3;
    end
    if (reset) begin
      reg_B_3_1_4 <= 32'sh0;
    end else begin
      reg_B_3_1_4 <= io_in_B_5_4;
    end
    if (reset) begin
      reg_B_3_1_5 <= 32'sh0;
    end else begin
      reg_B_3_1_5 <= io_in_B_5_5;
    end
    if (reset) begin
      reg_B_3_1_6 <= 32'sh0;
    end else begin
      reg_B_3_1_6 <= io_in_B_5_6;
    end
    if (reset) begin
      reg_B_3_1_7 <= 32'sh0;
    end else begin
      reg_B_3_1_7 <= io_in_B_5_7;
    end
    if (reset) begin
      reg_B_3_2_0 <= 32'sh0;
    end else begin
      reg_B_3_2_0 <= io_in_B_6_0;
    end
    if (reset) begin
      reg_B_3_2_1 <= 32'sh0;
    end else begin
      reg_B_3_2_1 <= io_in_B_6_1;
    end
    if (reset) begin
      reg_B_3_2_2 <= 32'sh0;
    end else begin
      reg_B_3_2_2 <= io_in_B_6_2;
    end
    if (reset) begin
      reg_B_3_2_3 <= 32'sh0;
    end else begin
      reg_B_3_2_3 <= io_in_B_6_3;
    end
    if (reset) begin
      reg_B_3_2_4 <= 32'sh0;
    end else begin
      reg_B_3_2_4 <= io_in_B_6_4;
    end
    if (reset) begin
      reg_B_3_2_5 <= 32'sh0;
    end else begin
      reg_B_3_2_5 <= io_in_B_6_5;
    end
    if (reset) begin
      reg_B_3_2_6 <= 32'sh0;
    end else begin
      reg_B_3_2_6 <= io_in_B_6_6;
    end
    if (reset) begin
      reg_B_3_2_7 <= 32'sh0;
    end else begin
      reg_B_3_2_7 <= io_in_B_6_7;
    end
    if (reset) begin
      reg_B_3_3_0 <= 32'sh0;
    end else begin
      reg_B_3_3_0 <= io_in_B_7_0;
    end
    if (reset) begin
      reg_B_3_3_1 <= 32'sh0;
    end else begin
      reg_B_3_3_1 <= io_in_B_7_1;
    end
    if (reset) begin
      reg_B_3_3_2 <= 32'sh0;
    end else begin
      reg_B_3_3_2 <= io_in_B_7_2;
    end
    if (reset) begin
      reg_B_3_3_3 <= 32'sh0;
    end else begin
      reg_B_3_3_3 <= io_in_B_7_3;
    end
    if (reset) begin
      reg_B_3_3_4 <= 32'sh0;
    end else begin
      reg_B_3_3_4 <= io_in_B_7_4;
    end
    if (reset) begin
      reg_B_3_3_5 <= 32'sh0;
    end else begin
      reg_B_3_3_5 <= io_in_B_7_5;
    end
    if (reset) begin
      reg_B_3_3_6 <= 32'sh0;
    end else begin
      reg_B_3_3_6 <= io_in_B_7_6;
    end
    if (reset) begin
      reg_B_3_3_7 <= 32'sh0;
    end else begin
      reg_B_3_3_7 <= io_in_B_7_7;
    end
    if (reset) begin
      reg_B_4_0_0 <= 32'sh0;
    end else begin
      reg_B_4_0_0 <= io_in_B_4_8;
    end
    if (reset) begin
      reg_B_4_0_1 <= 32'sh0;
    end else begin
      reg_B_4_0_1 <= io_in_B_4_9;
    end
    if (reset) begin
      reg_B_4_0_2 <= 32'sh0;
    end else begin
      reg_B_4_0_2 <= io_in_B_4_10;
    end
    if (reset) begin
      reg_B_4_0_3 <= 32'sh0;
    end else begin
      reg_B_4_0_3 <= io_in_B_4_11;
    end
    if (reset) begin
      reg_B_4_0_4 <= 32'sh0;
    end else begin
      reg_B_4_0_4 <= io_in_B_4_12;
    end
    if (reset) begin
      reg_B_4_0_5 <= 32'sh0;
    end else begin
      reg_B_4_0_5 <= io_in_B_4_13;
    end
    if (reset) begin
      reg_B_4_0_6 <= 32'sh0;
    end else begin
      reg_B_4_0_6 <= io_in_B_4_14;
    end
    if (reset) begin
      reg_B_4_0_7 <= 32'sh0;
    end else begin
      reg_B_4_0_7 <= io_in_B_4_15;
    end
    if (reset) begin
      reg_B_4_1_0 <= 32'sh0;
    end else begin
      reg_B_4_1_0 <= io_in_B_5_8;
    end
    if (reset) begin
      reg_B_4_1_1 <= 32'sh0;
    end else begin
      reg_B_4_1_1 <= io_in_B_5_9;
    end
    if (reset) begin
      reg_B_4_1_2 <= 32'sh0;
    end else begin
      reg_B_4_1_2 <= io_in_B_5_10;
    end
    if (reset) begin
      reg_B_4_1_3 <= 32'sh0;
    end else begin
      reg_B_4_1_3 <= io_in_B_5_11;
    end
    if (reset) begin
      reg_B_4_1_4 <= 32'sh0;
    end else begin
      reg_B_4_1_4 <= io_in_B_5_12;
    end
    if (reset) begin
      reg_B_4_1_5 <= 32'sh0;
    end else begin
      reg_B_4_1_5 <= io_in_B_5_13;
    end
    if (reset) begin
      reg_B_4_1_6 <= 32'sh0;
    end else begin
      reg_B_4_1_6 <= io_in_B_5_14;
    end
    if (reset) begin
      reg_B_4_1_7 <= 32'sh0;
    end else begin
      reg_B_4_1_7 <= io_in_B_5_15;
    end
    if (reset) begin
      reg_B_4_2_0 <= 32'sh0;
    end else begin
      reg_B_4_2_0 <= io_in_B_6_8;
    end
    if (reset) begin
      reg_B_4_2_1 <= 32'sh0;
    end else begin
      reg_B_4_2_1 <= io_in_B_6_9;
    end
    if (reset) begin
      reg_B_4_2_2 <= 32'sh0;
    end else begin
      reg_B_4_2_2 <= io_in_B_6_10;
    end
    if (reset) begin
      reg_B_4_2_3 <= 32'sh0;
    end else begin
      reg_B_4_2_3 <= io_in_B_6_11;
    end
    if (reset) begin
      reg_B_4_2_4 <= 32'sh0;
    end else begin
      reg_B_4_2_4 <= io_in_B_6_12;
    end
    if (reset) begin
      reg_B_4_2_5 <= 32'sh0;
    end else begin
      reg_B_4_2_5 <= io_in_B_6_13;
    end
    if (reset) begin
      reg_B_4_2_6 <= 32'sh0;
    end else begin
      reg_B_4_2_6 <= io_in_B_6_14;
    end
    if (reset) begin
      reg_B_4_2_7 <= 32'sh0;
    end else begin
      reg_B_4_2_7 <= io_in_B_6_15;
    end
    if (reset) begin
      reg_B_4_3_0 <= 32'sh0;
    end else begin
      reg_B_4_3_0 <= io_in_B_7_8;
    end
    if (reset) begin
      reg_B_4_3_1 <= 32'sh0;
    end else begin
      reg_B_4_3_1 <= io_in_B_7_9;
    end
    if (reset) begin
      reg_B_4_3_2 <= 32'sh0;
    end else begin
      reg_B_4_3_2 <= io_in_B_7_10;
    end
    if (reset) begin
      reg_B_4_3_3 <= 32'sh0;
    end else begin
      reg_B_4_3_3 <= io_in_B_7_11;
    end
    if (reset) begin
      reg_B_4_3_4 <= 32'sh0;
    end else begin
      reg_B_4_3_4 <= io_in_B_7_12;
    end
    if (reset) begin
      reg_B_4_3_5 <= 32'sh0;
    end else begin
      reg_B_4_3_5 <= io_in_B_7_13;
    end
    if (reset) begin
      reg_B_4_3_6 <= 32'sh0;
    end else begin
      reg_B_4_3_6 <= io_in_B_7_14;
    end
    if (reset) begin
      reg_B_4_3_7 <= 32'sh0;
    end else begin
      reg_B_4_3_7 <= io_in_B_7_15;
    end
    if (reset) begin
      cal_state_0 <= 1'h0;
    end else begin
      cal_state_0 <= TPUs_0_out_cal;
    end
    if (reset) begin
      cal_state_1 <= 1'h0;
    end else begin
      cal_state_1 <= _T_40965;
    end
    if (reset) begin
      cal_state_2 <= 1'h0;
    end else begin
      cal_state_2 <= TPUs_3_out_cal;
    end
    if (reset) begin
      result_0_0 <= 32'sh0;
    end else begin
      result_0_0 <= TPUs_0_out_result_0_0;
    end
    if (reset) begin
      result_0_1 <= 32'sh0;
    end else begin
      result_0_1 <= TPUs_0_out_result_0_1;
    end
    if (reset) begin
      result_0_2 <= 32'sh0;
    end else begin
      result_0_2 <= TPUs_0_out_result_0_2;
    end
    if (reset) begin
      result_0_3 <= 32'sh0;
    end else begin
      result_0_3 <= TPUs_0_out_result_0_3;
    end
    if (reset) begin
      result_0_4 <= 32'sh0;
    end else begin
      result_0_4 <= TPUs_1_out_result_0_0;
    end
    if (reset) begin
      result_0_5 <= 32'sh0;
    end else begin
      result_0_5 <= TPUs_1_out_result_0_1;
    end
    if (reset) begin
      result_0_6 <= 32'sh0;
    end else begin
      result_0_6 <= TPUs_1_out_result_0_2;
    end
    if (reset) begin
      result_0_7 <= 32'sh0;
    end else begin
      result_0_7 <= TPUs_1_out_result_0_3;
    end
    if (reset) begin
      result_1_0 <= 32'sh0;
    end else begin
      result_1_0 <= TPUs_0_out_result_1_0;
    end
    if (reset) begin
      result_1_1 <= 32'sh0;
    end else begin
      result_1_1 <= TPUs_0_out_result_1_1;
    end
    if (reset) begin
      result_1_2 <= 32'sh0;
    end else begin
      result_1_2 <= TPUs_0_out_result_1_2;
    end
    if (reset) begin
      result_1_3 <= 32'sh0;
    end else begin
      result_1_3 <= TPUs_0_out_result_1_3;
    end
    if (reset) begin
      result_1_4 <= 32'sh0;
    end else begin
      result_1_4 <= TPUs_1_out_result_1_0;
    end
    if (reset) begin
      result_1_5 <= 32'sh0;
    end else begin
      result_1_5 <= TPUs_1_out_result_1_1;
    end
    if (reset) begin
      result_1_6 <= 32'sh0;
    end else begin
      result_1_6 <= TPUs_1_out_result_1_2;
    end
    if (reset) begin
      result_1_7 <= 32'sh0;
    end else begin
      result_1_7 <= TPUs_1_out_result_1_3;
    end
    if (reset) begin
      result_2_0 <= 32'sh0;
    end else begin
      result_2_0 <= TPUs_2_out_result_0_0;
    end
    if (reset) begin
      result_2_1 <= 32'sh0;
    end else begin
      result_2_1 <= TPUs_2_out_result_0_1;
    end
    if (reset) begin
      result_2_2 <= 32'sh0;
    end else begin
      result_2_2 <= TPUs_2_out_result_0_2;
    end
    if (reset) begin
      result_2_3 <= 32'sh0;
    end else begin
      result_2_3 <= TPUs_2_out_result_0_3;
    end
    if (reset) begin
      result_2_4 <= 32'sh0;
    end else begin
      result_2_4 <= TPUs_3_out_result_0_0;
    end
    if (reset) begin
      result_2_5 <= 32'sh0;
    end else begin
      result_2_5 <= TPUs_3_out_result_0_1;
    end
    if (reset) begin
      result_2_6 <= 32'sh0;
    end else begin
      result_2_6 <= TPUs_3_out_result_0_2;
    end
    if (reset) begin
      result_2_7 <= 32'sh0;
    end else begin
      result_2_7 <= TPUs_3_out_result_0_3;
    end
    if (reset) begin
      result_3_0 <= 32'sh0;
    end else begin
      result_3_0 <= TPUs_2_out_result_1_0;
    end
    if (reset) begin
      result_3_1 <= 32'sh0;
    end else begin
      result_3_1 <= TPUs_2_out_result_1_1;
    end
    if (reset) begin
      result_3_2 <= 32'sh0;
    end else begin
      result_3_2 <= TPUs_2_out_result_1_2;
    end
    if (reset) begin
      result_3_3 <= 32'sh0;
    end else begin
      result_3_3 <= TPUs_2_out_result_1_3;
    end
    if (reset) begin
      result_3_4 <= 32'sh0;
    end else begin
      result_3_4 <= TPUs_3_out_result_1_0;
    end
    if (reset) begin
      result_3_5 <= 32'sh0;
    end else begin
      result_3_5 <= TPUs_3_out_result_1_1;
    end
    if (reset) begin
      result_3_6 <= 32'sh0;
    end else begin
      result_3_6 <= TPUs_3_out_result_1_2;
    end
    if (reset) begin
      result_3_7 <= 32'sh0;
    end else begin
      result_3_7 <= TPUs_3_out_result_1_3;
    end
    if (reset) begin
      cal_control_0 <= 1'h0;
    end else begin
      if (!(_T_43000)) begin
        if (_T_43006) begin
          if (!(_T_43007)) begin
            if (loop_reg) begin
              if (cal_state_0) begin
                cal_control_0 <= 1'h0;
              end else begin
                cal_control_0 <= 1'h1;
              end
            end
          end
        end else begin
          if (!(_T_43011)) begin
            if (_T_43016) begin
              if (!(_T_43007)) begin
                if (loop_reg) begin
                  if (_T_43021) begin
                    cal_control_0 <= 1'h0;
                  end else begin
                    cal_control_0 <= 1'h1;
                  end
                end
              end
            end else begin
              if (!(_T_43024)) begin
                if (_T_43029) begin
                  if (!(_T_43007)) begin
                    if (loop_reg) begin
                      if (cal_state_2) begin
                        cal_control_0 <= 1'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cal_control_1 <= 1'h0;
    end else begin
      if (!(_T_43000)) begin
        if (!(_T_43006)) begin
          if (_T_43011) begin
            if (!(_T_43007)) begin
              if (loop_reg) begin
                if (cal_state_1) begin
                  cal_control_1 <= 1'h0;
                end else begin
                  cal_control_1 <= 1'h1;
                end
              end
            end
          end else begin
            if (!(_T_43016)) begin
              if (_T_43024) begin
                if (!(_T_43007)) begin
                  if (loop_reg) begin
                    if (cal_state_1) begin
                      cal_control_1 <= 1'h0;
                    end else begin
                      cal_control_1 <= 1'h1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      cal_control_2 <= 1'h0;
    end else begin
      if (!(_T_43000)) begin
        if (!(_T_43006)) begin
          if (!(_T_43011)) begin
            if (_T_43016) begin
              if (!(_T_43007)) begin
                if (loop_reg) begin
                  if (_T_43021) begin
                    cal_control_2 <= 1'h0;
                  end else begin
                    cal_control_2 <= 1'h1;
                  end
                end
              end
            end else begin
              if (!(_T_43024)) begin
                if (_T_43029) begin
                  if (!(_T_43007)) begin
                    if (loop_reg) begin
                      cal_control_2 <= 1'h1;
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      stateReg <= 3'h0;
    end else begin
      if (_T_43000) begin
        if (_T_43005) begin
          stateReg <= 3'h1;
        end
      end else begin
        if (_T_43006) begin
          if (!(_T_43007)) begin
            if (loop_reg) begin
              if (cal_state_0) begin
                stateReg <= 3'h2;
              end
            end
          end
        end else begin
          if (_T_43011) begin
            if (!(_T_43007)) begin
              if (loop_reg) begin
                if (cal_state_1) begin
                  stateReg <= 3'h3;
                end
              end
            end
          end else begin
            if (_T_43016) begin
              if (!(_T_43007)) begin
                if (loop_reg) begin
                  if (_T_43021) begin
                    stateReg <= 3'h4;
                  end
                end
              end
            end else begin
              if (_T_43024) begin
                if (!(_T_43007)) begin
                  if (loop_reg) begin
                    if (cal_state_1) begin
                      stateReg <= 3'h5;
                    end
                  end
                end
              end else begin
                if (_T_43029) begin
                  if (!(_T_43007)) begin
                    if (loop_reg) begin
                      if (cal_state_2) begin
                        stateReg <= 3'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    if (reset) begin
      loop_reg <= 1'h0;
    end else begin
      if (!(_T_43000)) begin
        if (_T_43006) begin
          if (_T_43007) begin
            loop_reg <= 1'h1;
          end else begin
            if (loop_reg) begin
              if (cal_state_0) begin
                loop_reg <= 1'h0;
              end
            end
          end
        end else begin
          if (_T_43011) begin
            if (_T_43007) begin
              loop_reg <= 1'h1;
            end else begin
              if (loop_reg) begin
                if (cal_state_1) begin
                  loop_reg <= 1'h0;
                end
              end
            end
          end else begin
            if (_T_43016) begin
              if (_T_43007) begin
                loop_reg <= 1'h1;
              end else begin
                if (loop_reg) begin
                  if (_T_43021) begin
                    loop_reg <= 1'h0;
                  end
                end
              end
            end else begin
              if (_T_43024) begin
                if (_T_43007) begin
                  loop_reg <= 1'h1;
                end else begin
                  if (loop_reg) begin
                    if (cal_state_1) begin
                      loop_reg <= 1'h0;
                    end
                  end
                end
              end else begin
                if (_T_43029) begin
                  if (_T_43007) begin
                    loop_reg <= 1'h1;
                  end else begin
                    if (loop_reg) begin
                      if (cal_state_2) begin
                        loop_reg <= 1'h0;
                      end
                    end
                  end
                end
              end
            end
          end
        end
      end
    end
    _T_43002 <= io_in_cal;
  end
endmodule
