module tag( // @[:@3.2]
  input clock, // @[:@4.4]
  input reset, // @[:@5.4]
  output io_out_tag_0, // @[:@6.4]
  output io_out_tag_1, // @[:@6.4]
  output io_out_tag_2, // @[:@6.4]
  output io_out_tag_3, // @[:@6.4]
  output io_out_tag_4, // @[:@6.4]
  output io_out_tag_5, // @[:@6.4]
  output io_out_tag_6 // @[:@6.4]
);
  reg tag_0; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_0;
  reg tag_1; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_1;
  reg tag_2; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_2;
  reg tag_3; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_3;
  reg tag_4; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_4;
  reg tag_5; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_5;
  reg tag_6; // @[tag.scala 32:20:@17.4]
  reg [31:0] _RAND_6;
  assign io_out_tag_0 = tag_0; // @[tag.scala 42:14:@47.4]
  assign io_out_tag_1 = tag_1; // @[tag.scala 42:14:@48.4]
  assign io_out_tag_2 = tag_2; // @[tag.scala 42:14:@49.4]
  assign io_out_tag_3 = tag_3; // @[tag.scala 42:14:@50.4]
  assign io_out_tag_4 = tag_4; // @[tag.scala 42:14:@51.4]
  assign io_out_tag_5 = tag_5; // @[tag.scala 42:14:@52.4]
  assign io_out_tag_6 = tag_6; // @[tag.scala 42:14:@53.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  tag_0 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  tag_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  tag_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  tag_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  tag_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  tag_5 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  tag_6 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      tag_0 <= 1'h0;
    end else begin
      tag_0 <= 1'h1;
    end
    if (reset) begin
      tag_1 <= 1'h0;
    end else begin
      tag_1 <= 1'h1;
    end
    if (reset) begin
      tag_2 <= 1'h0;
    end else begin
      tag_2 <= 1'h1;
    end
    if (reset) begin
      tag_3 <= 1'h0;
    end else begin
      tag_3 <= 1'h1;
    end
    if (reset) begin
      tag_4 <= 1'h0;
    end else begin
      tag_4 <= 1'h1;
    end
    if (reset) begin
      tag_5 <= 1'h0;
    end else begin
      tag_5 <= 1'h1;
    end
    if (reset) begin
      tag_6 <= 1'h0;
    end else begin
      tag_6 <= 1'h1;
    end
  end
endmodule
module MUX8( // @[:@219.2]
  input [31:0] io_int_in_0, // @[:@222.4]
  input [31:0] io_int_in_1, // @[:@222.4]
  input [31:0] io_int_in_2, // @[:@222.4]
  input [31:0] io_int_in_3, // @[:@222.4]
  input [31:0] io_int_in_4, // @[:@222.4]
  input [31:0] io_int_in_5, // @[:@222.4]
  input [31:0] io_int_in_6, // @[:@222.4]
  input [31:0] io_int_in_7, // @[:@222.4]
  input io_tag_0, // @[:@222.4]
  input io_tag_1, // @[:@222.4]
  input io_tag_2, // @[:@222.4]
  input io_tag_3, // @[:@222.4]
  input io_tag_4, // @[:@222.4]
  input io_tag_5, // @[:@222.4]
  input io_tag_6, // @[:@222.4]
  input io_tag_7, // @[:@222.4]
  output [31:0] io_choice // @[:@222.4]
);
  wire [31:0] _T_62; // @[Mux.scala 19:72:@225.4]
  wire [31:0] _T_63; // @[Mux.scala 19:72:@226.4]
  wire [31:0] _T_66; // @[Mux.scala 19:72:@229.4]
  wire [31:0] _T_67; // @[Mux.scala 19:72:@230.4]
  wire [31:0] _T_70; // @[Mux.scala 19:72:@233.4]
  wire [31:0] _T_71; // @[Mux.scala 19:72:@234.4]
  wire [31:0] _T_74; // @[Mux.scala 19:72:@237.4]
  wire [31:0] _T_75; // @[Mux.scala 19:72:@238.4]
  wire [31:0] _T_78; // @[Mux.scala 19:72:@241.4]
  wire [31:0] _T_79; // @[Mux.scala 19:72:@242.4]
  wire [31:0] _T_82; // @[Mux.scala 19:72:@245.4]
  wire [31:0] _T_83; // @[Mux.scala 19:72:@246.4]
  wire [31:0] _T_86; // @[Mux.scala 19:72:@249.4]
  wire [31:0] _T_87; // @[Mux.scala 19:72:@250.4]
  wire [31:0] _T_90; // @[Mux.scala 19:72:@253.4]
  wire [31:0] _T_91; // @[Mux.scala 19:72:@254.4]
  wire [31:0] _T_93; // @[Mux.scala 19:72:@256.4]
  wire [31:0] _T_95; // @[Mux.scala 19:72:@257.4]
  wire [31:0] _T_97; // @[Mux.scala 19:72:@258.4]
  wire [31:0] _T_99; // @[Mux.scala 19:72:@259.4]
  wire [31:0] _T_101; // @[Mux.scala 19:72:@260.4]
  wire [31:0] _T_103; // @[Mux.scala 19:72:@261.4]
  wire [31:0] _T_105; // @[Mux.scala 19:72:@262.4]
  wire [31:0] _T_107; // @[Mux.scala 19:72:@263.4]
  wire [31:0] _T_108; // @[Mux.scala 19:72:@264.4]
  wire [31:0] _T_109; // @[Mux.scala 19:72:@265.4]
  wire [31:0] _T_110; // @[Mux.scala 19:72:@266.4]
  wire [31:0] _T_111; // @[Mux.scala 19:72:@267.4]
  wire [31:0] _T_112; // @[Mux.scala 19:72:@268.4]
  wire [31:0] _T_113; // @[Mux.scala 19:72:@269.4]
  wire [31:0] _T_114; // @[Mux.scala 19:72:@270.4]
  wire [31:0] _T_115; // @[Mux.scala 19:72:@271.4]
  wire [31:0] _T_116; // @[Mux.scala 19:72:@272.4]
  wire [31:0] _T_117; // @[Mux.scala 19:72:@273.4]
  wire [31:0] _T_118; // @[Mux.scala 19:72:@274.4]
  wire [31:0] _T_119; // @[Mux.scala 19:72:@275.4]
  wire [31:0] _T_120; // @[Mux.scala 19:72:@276.4]
  wire [31:0] _T_121; // @[Mux.scala 19:72:@277.4]
  wire [31:0] _T_124; // @[Mux.scala 19:72:@279.4]
  assign _T_62 = $unsigned(io_int_in_0); // @[Mux.scala 19:72:@225.4]
  assign _T_63 = $signed(_T_62); // @[Mux.scala 19:72:@226.4]
  assign _T_66 = $unsigned(io_int_in_1); // @[Mux.scala 19:72:@229.4]
  assign _T_67 = $signed(_T_66); // @[Mux.scala 19:72:@230.4]
  assign _T_70 = $unsigned(io_int_in_2); // @[Mux.scala 19:72:@233.4]
  assign _T_71 = $signed(_T_70); // @[Mux.scala 19:72:@234.4]
  assign _T_74 = $unsigned(io_int_in_3); // @[Mux.scala 19:72:@237.4]
  assign _T_75 = $signed(_T_74); // @[Mux.scala 19:72:@238.4]
  assign _T_78 = $unsigned(io_int_in_4); // @[Mux.scala 19:72:@241.4]
  assign _T_79 = $signed(_T_78); // @[Mux.scala 19:72:@242.4]
  assign _T_82 = $unsigned(io_int_in_5); // @[Mux.scala 19:72:@245.4]
  assign _T_83 = $signed(_T_82); // @[Mux.scala 19:72:@246.4]
  assign _T_86 = $unsigned(io_int_in_6); // @[Mux.scala 19:72:@249.4]
  assign _T_87 = $signed(_T_86); // @[Mux.scala 19:72:@250.4]
  assign _T_90 = $unsigned(io_int_in_7); // @[Mux.scala 19:72:@253.4]
  assign _T_91 = $signed(_T_90); // @[Mux.scala 19:72:@254.4]
  assign _T_93 = io_tag_0 ? $signed(_T_63):$signed(32'sh0); // @[Mux.scala 19:72:@256.4]
  assign _T_95 = io_tag_1 ? $signed(_T_67):$signed(32'sh0); // @[Mux.scala 19:72:@257.4]
  assign _T_97 = io_tag_2 ? $signed(_T_71):$signed(32'sh0); // @[Mux.scala 19:72:@258.4]
  assign _T_99 = io_tag_3 ? $signed(_T_75):$signed(32'sh0); // @[Mux.scala 19:72:@259.4]
  assign _T_101 = io_tag_4 ? $signed(_T_79):$signed(32'sh0); // @[Mux.scala 19:72:@260.4]
  assign _T_103 = io_tag_5 ? $signed(_T_83):$signed(32'sh0); // @[Mux.scala 19:72:@261.4]
  assign _T_105 = io_tag_6 ? $signed(_T_87):$signed(32'sh0); // @[Mux.scala 19:72:@262.4]
  assign _T_107 = io_tag_7 ? $signed(_T_91):$signed(32'sh0); // @[Mux.scala 19:72:@263.4]
  assign _T_108 = $signed(_T_93) | $signed(_T_95); // @[Mux.scala 19:72:@264.4]
  assign _T_109 = $signed(_T_108); // @[Mux.scala 19:72:@265.4]
  assign _T_110 = $signed(_T_109) | $signed(_T_97); // @[Mux.scala 19:72:@266.4]
  assign _T_111 = $signed(_T_110); // @[Mux.scala 19:72:@267.4]
  assign _T_112 = $signed(_T_111) | $signed(_T_99); // @[Mux.scala 19:72:@268.4]
  assign _T_113 = $signed(_T_112); // @[Mux.scala 19:72:@269.4]
  assign _T_114 = $signed(_T_113) | $signed(_T_101); // @[Mux.scala 19:72:@270.4]
  assign _T_115 = $signed(_T_114); // @[Mux.scala 19:72:@271.4]
  assign _T_116 = $signed(_T_115) | $signed(_T_103); // @[Mux.scala 19:72:@272.4]
  assign _T_117 = $signed(_T_116); // @[Mux.scala 19:72:@273.4]
  assign _T_118 = $signed(_T_117) | $signed(_T_105); // @[Mux.scala 19:72:@274.4]
  assign _T_119 = $signed(_T_118); // @[Mux.scala 19:72:@275.4]
  assign _T_120 = $signed(_T_119) | $signed(_T_107); // @[Mux.scala 19:72:@276.4]
  assign _T_121 = $signed(_T_120); // @[Mux.scala 19:72:@277.4]
  assign _T_124 = $unsigned(_T_121); // @[Mux.scala 19:72:@279.4]
  assign io_choice = $signed(_T_124); // @[MUX8.scala 40:13:@282.4]
endmodule
module tag_refine( // @[:@544.2]
  input clock, // @[:@545.4]
  input reset, // @[:@546.4]
  input io_tag_in_0, // @[:@547.4]
  input io_tag_in_1, // @[:@547.4]
  input io_tag_in_2, // @[:@547.4]
  input io_tag_in_3, // @[:@547.4]
  input io_tag_in_4, // @[:@547.4]
  input io_tag_in_5, // @[:@547.4]
  input io_tag_in_6, // @[:@547.4]
  input io_tag_in_7, // @[:@547.4]
  output io_tag_out_0, // @[:@547.4]
  output io_tag_out_1, // @[:@547.4]
  output io_tag_out_2, // @[:@547.4]
  output io_tag_out_3, // @[:@547.4]
  output io_tag_out_4, // @[:@547.4]
  output io_tag_out_5, // @[:@547.4]
  output io_tag_out_6, // @[:@547.4]
  output io_tag_out_7 // @[:@547.4]
);
  reg tag_0; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_0;
  reg tag_1; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_1;
  reg tag_2; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_2;
  reg tag_3; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_3;
  reg tag_4; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_4;
  reg tag_5; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_5;
  reg tag_6; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_6;
  reg tag_7; // @[tag_refine.scala 28:20:@558.4]
  reg [31:0] _RAND_7;
  reg find; // @[tag_refine.scala 29:21:@559.4]
  reg [31:0] _RAND_8;
  wire _T_130; // @[tag_refine.scala 34:15:@568.4]
  wire _GEN_0; // @[tag_refine.scala 35:31:@571.6]
  wire _GEN_1; // @[tag_refine.scala 35:31:@571.6]
  wire _GEN_2; // @[tag_refine.scala 34:28:@569.4]
  wire _GEN_3; // @[tag_refine.scala 34:28:@569.4]
  wire _GEN_4; // @[tag_refine.scala 35:31:@579.6]
  wire _GEN_5; // @[tag_refine.scala 35:31:@579.6]
  wire _GEN_6; // @[tag_refine.scala 34:28:@577.4]
  wire _GEN_7; // @[tag_refine.scala 34:28:@577.4]
  wire _GEN_8; // @[tag_refine.scala 35:31:@587.6]
  wire _GEN_9; // @[tag_refine.scala 35:31:@587.6]
  wire _GEN_10; // @[tag_refine.scala 34:28:@585.4]
  wire _GEN_11; // @[tag_refine.scala 34:28:@585.4]
  wire _GEN_12; // @[tag_refine.scala 35:31:@595.6]
  wire _GEN_13; // @[tag_refine.scala 35:31:@595.6]
  wire _GEN_14; // @[tag_refine.scala 34:28:@593.4]
  wire _GEN_15; // @[tag_refine.scala 34:28:@593.4]
  wire _GEN_16; // @[tag_refine.scala 35:31:@603.6]
  wire _GEN_17; // @[tag_refine.scala 35:31:@603.6]
  wire _GEN_18; // @[tag_refine.scala 34:28:@601.4]
  wire _GEN_19; // @[tag_refine.scala 34:28:@601.4]
  wire _GEN_20; // @[tag_refine.scala 35:31:@611.6]
  wire _GEN_21; // @[tag_refine.scala 35:31:@611.6]
  wire _GEN_22; // @[tag_refine.scala 34:28:@609.4]
  wire _GEN_23; // @[tag_refine.scala 34:28:@609.4]
  wire _GEN_24; // @[tag_refine.scala 35:31:@619.6]
  wire _GEN_25; // @[tag_refine.scala 35:31:@619.6]
  wire _GEN_26; // @[tag_refine.scala 34:28:@617.4]
  wire _GEN_27; // @[tag_refine.scala 34:28:@617.4]
  wire _GEN_28; // @[tag_refine.scala 35:31:@627.6]
  wire _GEN_29; // @[tag_refine.scala 35:31:@627.6]
  wire _GEN_30; // @[tag_refine.scala 34:28:@625.4]
  wire _GEN_31; // @[tag_refine.scala 34:28:@625.4]
  assign _T_130 = find == 1'h0; // @[tag_refine.scala 34:15:@568.4]
  assign _GEN_0 = tag_0 ? 1'h0:io_tag_in_0; // @[tag_refine.scala 35:31:@571.6]
  assign _GEN_1 = tag_0 ? 1'h1:find; // @[tag_refine.scala 35:31:@571.6]
  assign _GEN_2 = _T_130 ? _GEN_0:io_tag_in_0; // @[tag_refine.scala 34:28:@569.4]
  assign _GEN_3 = _T_130 ? _GEN_1:find; // @[tag_refine.scala 34:28:@569.4]
  assign _GEN_4 = tag_1 ? 1'h0:io_tag_in_1; // @[tag_refine.scala 35:31:@579.6]
  assign _GEN_5 = tag_1 ? 1'h1:_GEN_3; // @[tag_refine.scala 35:31:@579.6]
  assign _GEN_6 = _T_130 ? _GEN_4:io_tag_in_1; // @[tag_refine.scala 34:28:@577.4]
  assign _GEN_7 = _T_130 ? _GEN_5:_GEN_3; // @[tag_refine.scala 34:28:@577.4]
  assign _GEN_8 = tag_2 ? 1'h0:io_tag_in_2; // @[tag_refine.scala 35:31:@587.6]
  assign _GEN_9 = tag_2 ? 1'h1:_GEN_7; // @[tag_refine.scala 35:31:@587.6]
  assign _GEN_10 = _T_130 ? _GEN_8:io_tag_in_2; // @[tag_refine.scala 34:28:@585.4]
  assign _GEN_11 = _T_130 ? _GEN_9:_GEN_7; // @[tag_refine.scala 34:28:@585.4]
  assign _GEN_12 = tag_3 ? 1'h0:io_tag_in_3; // @[tag_refine.scala 35:31:@595.6]
  assign _GEN_13 = tag_3 ? 1'h1:_GEN_11; // @[tag_refine.scala 35:31:@595.6]
  assign _GEN_14 = _T_130 ? _GEN_12:io_tag_in_3; // @[tag_refine.scala 34:28:@593.4]
  assign _GEN_15 = _T_130 ? _GEN_13:_GEN_11; // @[tag_refine.scala 34:28:@593.4]
  assign _GEN_16 = tag_4 ? 1'h0:io_tag_in_4; // @[tag_refine.scala 35:31:@603.6]
  assign _GEN_17 = tag_4 ? 1'h1:_GEN_15; // @[tag_refine.scala 35:31:@603.6]
  assign _GEN_18 = _T_130 ? _GEN_16:io_tag_in_4; // @[tag_refine.scala 34:28:@601.4]
  assign _GEN_19 = _T_130 ? _GEN_17:_GEN_15; // @[tag_refine.scala 34:28:@601.4]
  assign _GEN_20 = tag_5 ? 1'h0:io_tag_in_5; // @[tag_refine.scala 35:31:@611.6]
  assign _GEN_21 = tag_5 ? 1'h1:_GEN_19; // @[tag_refine.scala 35:31:@611.6]
  assign _GEN_22 = _T_130 ? _GEN_20:io_tag_in_5; // @[tag_refine.scala 34:28:@609.4]
  assign _GEN_23 = _T_130 ? _GEN_21:_GEN_19; // @[tag_refine.scala 34:28:@609.4]
  assign _GEN_24 = tag_6 ? 1'h0:io_tag_in_6; // @[tag_refine.scala 35:31:@619.6]
  assign _GEN_25 = tag_6 ? 1'h1:_GEN_23; // @[tag_refine.scala 35:31:@619.6]
  assign _GEN_26 = _T_130 ? _GEN_24:io_tag_in_6; // @[tag_refine.scala 34:28:@617.4]
  assign _GEN_27 = _T_130 ? _GEN_25:_GEN_23; // @[tag_refine.scala 34:28:@617.4]
  assign _GEN_28 = tag_7 ? 1'h0:io_tag_in_7; // @[tag_refine.scala 35:31:@627.6]
  assign _GEN_29 = tag_7 ? 1'h1:_GEN_27; // @[tag_refine.scala 35:31:@627.6]
  assign _GEN_30 = _T_130 ? _GEN_28:io_tag_in_7; // @[tag_refine.scala 34:28:@625.4]
  assign _GEN_31 = _T_130 ? _GEN_29:_GEN_27; // @[tag_refine.scala 34:28:@625.4]
  assign io_tag_out_0 = tag_0; // @[tag_refine.scala 42:14:@632.4]
  assign io_tag_out_1 = tag_1; // @[tag_refine.scala 42:14:@633.4]
  assign io_tag_out_2 = tag_2; // @[tag_refine.scala 42:14:@634.4]
  assign io_tag_out_3 = tag_3; // @[tag_refine.scala 42:14:@635.4]
  assign io_tag_out_4 = tag_4; // @[tag_refine.scala 42:14:@636.4]
  assign io_tag_out_5 = tag_5; // @[tag_refine.scala 42:14:@637.4]
  assign io_tag_out_6 = tag_6; // @[tag_refine.scala 42:14:@638.4]
  assign io_tag_out_7 = tag_7; // @[tag_refine.scala 42:14:@639.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  tag_0 = _RAND_0[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  tag_1 = _RAND_1[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  tag_2 = _RAND_2[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  tag_3 = _RAND_3[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  tag_4 = _RAND_4[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  tag_5 = _RAND_5[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  tag_6 = _RAND_6[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  tag_7 = _RAND_7[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  find = _RAND_8[0:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      tag_0 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_0) begin
          tag_0 <= 1'h0;
        end else begin
          tag_0 <= io_tag_in_0;
        end
      end else begin
        tag_0 <= io_tag_in_0;
      end
    end
    if (reset) begin
      tag_1 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_1) begin
          tag_1 <= 1'h0;
        end else begin
          tag_1 <= io_tag_in_1;
        end
      end else begin
        tag_1 <= io_tag_in_1;
      end
    end
    if (reset) begin
      tag_2 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_2) begin
          tag_2 <= 1'h0;
        end else begin
          tag_2 <= io_tag_in_2;
        end
      end else begin
        tag_2 <= io_tag_in_2;
      end
    end
    if (reset) begin
      tag_3 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_3) begin
          tag_3 <= 1'h0;
        end else begin
          tag_3 <= io_tag_in_3;
        end
      end else begin
        tag_3 <= io_tag_in_3;
      end
    end
    if (reset) begin
      tag_4 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_4) begin
          tag_4 <= 1'h0;
        end else begin
          tag_4 <= io_tag_in_4;
        end
      end else begin
        tag_4 <= io_tag_in_4;
      end
    end
    if (reset) begin
      tag_5 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_5) begin
          tag_5 <= 1'h0;
        end else begin
          tag_5 <= io_tag_in_5;
        end
      end else begin
        tag_5 <= io_tag_in_5;
      end
    end
    if (reset) begin
      tag_6 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_6) begin
          tag_6 <= 1'h0;
        end else begin
          tag_6 <= io_tag_in_6;
        end
      end else begin
        tag_6 <= io_tag_in_6;
      end
    end
    if (reset) begin
      tag_7 <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_7) begin
          tag_7 <= 1'h0;
        end else begin
          tag_7 <= io_tag_in_7;
        end
      end else begin
        tag_7 <= io_tag_in_7;
      end
    end
    if (reset) begin
      find <= 1'h0;
    end else begin
      if (_T_130) begin
        if (tag_7) begin
          find <= 1'h1;
        end else begin
          if (_T_130) begin
            if (tag_6) begin
              find <= 1'h1;
            end else begin
              if (_T_130) begin
                if (tag_5) begin
                  find <= 1'h1;
                end else begin
                  if (_T_130) begin
                    if (tag_4) begin
                      find <= 1'h1;
                    end else begin
                      if (_T_130) begin
                        if (tag_3) begin
                          find <= 1'h1;
                        end else begin
                          if (_T_130) begin
                            if (tag_2) begin
                              find <= 1'h1;
                            end else begin
                              if (_T_130) begin
                                if (tag_1) begin
                                  find <= 1'h1;
                                end else begin
                                  if (_T_130) begin
                                    if (tag_0) begin
                                      find <= 1'h1;
                                    end
                                  end
                                end
                              end else begin
                                if (_T_130) begin
                                  if (tag_0) begin
                                    find <= 1'h1;
                                  end
                                end
                              end
                            end
                          end else begin
                            if (_T_130) begin
                              if (tag_1) begin
                                find <= 1'h1;
                              end else begin
                                if (_T_130) begin
                                  if (tag_0) begin
                                    find <= 1'h1;
                                  end
                                end
                              end
                            end else begin
                              if (_T_130) begin
                                if (tag_0) begin
                                  find <= 1'h1;
                                end
                              end
                            end
                          end
                        end
                      end else begin
                        if (_T_130) begin
                          if (tag_2) begin
                            find <= 1'h1;
                          end else begin
                            if (_T_130) begin
                              if (tag_1) begin
                                find <= 1'h1;
                              end else begin
                                find <= _GEN_3;
                              end
                            end else begin
                              find <= _GEN_3;
                            end
                          end
                        end else begin
                          if (_T_130) begin
                            if (tag_1) begin
                              find <= 1'h1;
                            end else begin
                              find <= _GEN_3;
                            end
                          end else begin
                            find <= _GEN_3;
                          end
                        end
                      end
                    end
                  end else begin
                    if (_T_130) begin
                      if (tag_3) begin
                        find <= 1'h1;
                      end else begin
                        if (_T_130) begin
                          if (tag_2) begin
                            find <= 1'h1;
                          end else begin
                            find <= _GEN_7;
                          end
                        end else begin
                          find <= _GEN_7;
                        end
                      end
                    end else begin
                      if (_T_130) begin
                        if (tag_2) begin
                          find <= 1'h1;
                        end else begin
                          find <= _GEN_7;
                        end
                      end else begin
                        find <= _GEN_7;
                      end
                    end
                  end
                end
              end else begin
                if (_T_130) begin
                  if (tag_4) begin
                    find <= 1'h1;
                  end else begin
                    if (_T_130) begin
                      if (tag_3) begin
                        find <= 1'h1;
                      end else begin
                        find <= _GEN_11;
                      end
                    end else begin
                      find <= _GEN_11;
                    end
                  end
                end else begin
                  if (_T_130) begin
                    if (tag_3) begin
                      find <= 1'h1;
                    end else begin
                      find <= _GEN_11;
                    end
                  end else begin
                    find <= _GEN_11;
                  end
                end
              end
            end
          end else begin
            if (_T_130) begin
              if (tag_5) begin
                find <= 1'h1;
              end else begin
                if (_T_130) begin
                  if (tag_4) begin
                    find <= 1'h1;
                  end else begin
                    find <= _GEN_15;
                  end
                end else begin
                  find <= _GEN_15;
                end
              end
            end else begin
              if (_T_130) begin
                if (tag_4) begin
                  find <= 1'h1;
                end else begin
                  find <= _GEN_15;
                end
              end else begin
                find <= _GEN_15;
              end
            end
          end
        end
      end else begin
        if (_T_130) begin
          if (tag_6) begin
            find <= 1'h1;
          end else begin
            if (_T_130) begin
              if (tag_5) begin
                find <= 1'h1;
              end else begin
                find <= _GEN_19;
              end
            end else begin
              find <= _GEN_19;
            end
          end
        end else begin
          if (_T_130) begin
            if (tag_5) begin
              find <= 1'h1;
            end else begin
              find <= _GEN_19;
            end
          end else begin
            find <= _GEN_19;
          end
        end
      end
    end
  end
endmodule
module S8DP1( // @[:@641.2]
  input clock, // @[:@642.4]
  input reset, // @[:@643.4]
  input [31:0] io_int_in_A_0, // @[:@644.4]
  input [31:0] io_int_in_A_1, // @[:@644.4]
  input [31:0] io_int_in_A_2, // @[:@644.4]
  input [31:0] io_int_in_A_3, // @[:@644.4]
  input [31:0] io_int_in_A_4, // @[:@644.4]
  input [31:0] io_int_in_A_5, // @[:@644.4]
  input [31:0] io_int_in_A_6, // @[:@644.4]
  input [31:0] io_int_in_A_7, // @[:@644.4]
  input [31:0] io_int_in_B, // @[:@644.4]
  input io_tag_0, // @[:@644.4]
  input io_tag_1, // @[:@644.4]
  input io_tag_2, // @[:@644.4]
  input io_tag_3, // @[:@644.4]
  input io_tag_4, // @[:@644.4]
  input io_tag_5, // @[:@644.4]
  input io_tag_6, // @[:@644.4]
  input io_tag_7, // @[:@644.4]
  output io_out_tag_0, // @[:@644.4]
  output io_out_tag_1, // @[:@644.4]
  output io_out_tag_2, // @[:@644.4]
  output io_out_tag_3, // @[:@644.4]
  output io_out_tag_4, // @[:@644.4]
  output io_out_tag_5, // @[:@644.4]
  output io_out_tag_6, // @[:@644.4]
  output io_out_tag_7, // @[:@644.4]
  output [31:0] io_result // @[:@644.4]
);
  wire [31:0] mux_io_int_in_0; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_1; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_2; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_3; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_4; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_5; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_6; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_int_in_7; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_0; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_1; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_2; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_3; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_4; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_5; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_6; // @[S8DP1.scala 29:19:@647.4]
  wire mux_io_tag_7; // @[S8DP1.scala 29:19:@647.4]
  wire [31:0] mux_io_choice; // @[S8DP1.scala 29:19:@647.4]
  wire tag_change_clock; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_reset; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_0; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_1; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_2; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_3; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_4; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_5; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_6; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_in_7; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_0; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_1; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_2; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_3; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_4; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_5; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_6; // @[S8DP1.scala 30:26:@650.4]
  wire tag_change_io_tag_out_7; // @[S8DP1.scala 30:26:@650.4]
  reg [31:0] acc; // @[S8DP1.scala 28:20:@646.4]
  reg [31:0] _RAND_0;
  wire [63:0] _T_89; // @[S8DP1.scala 35:28:@669.4]
  wire [63:0] _GEN_0; // @[S8DP1.scala 35:14:@670.4]
  wire [64:0] _T_90; // @[S8DP1.scala 35:14:@670.4]
  wire [63:0] _T_91; // @[S8DP1.scala 35:14:@671.4]
  wire [63:0] _T_92; // @[S8DP1.scala 35:14:@672.4]
  wire [31:0] _GEN_1; // @[S8DP1.scala 35:7:@673.4]
  MUX8 mux( // @[S8DP1.scala 29:19:@647.4]
    .io_int_in_0(mux_io_int_in_0),
    .io_int_in_1(mux_io_int_in_1),
    .io_int_in_2(mux_io_int_in_2),
    .io_int_in_3(mux_io_int_in_3),
    .io_int_in_4(mux_io_int_in_4),
    .io_int_in_5(mux_io_int_in_5),
    .io_int_in_6(mux_io_int_in_6),
    .io_int_in_7(mux_io_int_in_7),
    .io_tag_0(mux_io_tag_0),
    .io_tag_1(mux_io_tag_1),
    .io_tag_2(mux_io_tag_2),
    .io_tag_3(mux_io_tag_3),
    .io_tag_4(mux_io_tag_4),
    .io_tag_5(mux_io_tag_5),
    .io_tag_6(mux_io_tag_6),
    .io_tag_7(mux_io_tag_7),
    .io_choice(mux_io_choice)
  );
  tag_refine tag_change( // @[S8DP1.scala 30:26:@650.4]
    .clock(tag_change_clock),
    .reset(tag_change_reset),
    .io_tag_in_0(tag_change_io_tag_in_0),
    .io_tag_in_1(tag_change_io_tag_in_1),
    .io_tag_in_2(tag_change_io_tag_in_2),
    .io_tag_in_3(tag_change_io_tag_in_3),
    .io_tag_in_4(tag_change_io_tag_in_4),
    .io_tag_in_5(tag_change_io_tag_in_5),
    .io_tag_in_6(tag_change_io_tag_in_6),
    .io_tag_in_7(tag_change_io_tag_in_7),
    .io_tag_out_0(tag_change_io_tag_out_0),
    .io_tag_out_1(tag_change_io_tag_out_1),
    .io_tag_out_2(tag_change_io_tag_out_2),
    .io_tag_out_3(tag_change_io_tag_out_3),
    .io_tag_out_4(tag_change_io_tag_out_4),
    .io_tag_out_5(tag_change_io_tag_out_5),
    .io_tag_out_6(tag_change_io_tag_out_6),
    .io_tag_out_7(tag_change_io_tag_out_7)
  );
  assign _T_89 = $signed(io_int_in_B)*$signed(mux_io_choice); // @[S8DP1.scala 35:28:@669.4]
  assign _GEN_0 = {{32{acc[31]}}, acc}; // @[S8DP1.scala 35:14:@670.4]
  assign _T_90 = $signed(_GEN_0)+$signed(_T_89); // @[S8DP1.scala 35:14:@670.4]
  assign _T_91 = _T_90[63:0]; // @[S8DP1.scala 35:14:@671.4]
  assign _T_92 = $signed(_T_91); // @[S8DP1.scala 35:14:@672.4]
  assign io_out_tag_0 = tag_change_io_tag_out_0; // @[S8DP1.scala 38:14:@682.4]
  assign io_out_tag_1 = tag_change_io_tag_out_1; // @[S8DP1.scala 38:14:@683.4]
  assign io_out_tag_2 = tag_change_io_tag_out_2; // @[S8DP1.scala 38:14:@684.4]
  assign io_out_tag_3 = tag_change_io_tag_out_3; // @[S8DP1.scala 38:14:@685.4]
  assign io_out_tag_4 = tag_change_io_tag_out_4; // @[S8DP1.scala 38:14:@686.4]
  assign io_out_tag_5 = tag_change_io_tag_out_5; // @[S8DP1.scala 38:14:@687.4]
  assign io_out_tag_6 = tag_change_io_tag_out_6; // @[S8DP1.scala 38:14:@688.4]
  assign io_out_tag_7 = tag_change_io_tag_out_7; // @[S8DP1.scala 38:14:@689.4]
  assign io_result = acc; // @[S8DP1.scala 40:13:@690.4]
  assign _GEN_1 = _T_92[31:0]; // @[S8DP1.scala 35:7:@673.4]
  assign mux_io_int_in_0 = io_int_in_A_0; // @[S8DP1.scala 32:17:@653.4]
  assign mux_io_int_in_1 = io_int_in_A_1; // @[S8DP1.scala 32:17:@654.4]
  assign mux_io_int_in_2 = io_int_in_A_2; // @[S8DP1.scala 32:17:@655.4]
  assign mux_io_int_in_3 = io_int_in_A_3; // @[S8DP1.scala 32:17:@656.4]
  assign mux_io_int_in_4 = io_int_in_A_4; // @[S8DP1.scala 32:17:@657.4]
  assign mux_io_int_in_5 = io_int_in_A_5; // @[S8DP1.scala 32:17:@658.4]
  assign mux_io_int_in_6 = io_int_in_A_6; // @[S8DP1.scala 32:17:@659.4]
  assign mux_io_int_in_7 = io_int_in_A_7; // @[S8DP1.scala 32:17:@660.4]
  assign mux_io_tag_0 = io_tag_0; // @[S8DP1.scala 33:14:@661.4]
  assign mux_io_tag_1 = io_tag_1; // @[S8DP1.scala 33:14:@662.4]
  assign mux_io_tag_2 = io_tag_2; // @[S8DP1.scala 33:14:@663.4]
  assign mux_io_tag_3 = io_tag_3; // @[S8DP1.scala 33:14:@664.4]
  assign mux_io_tag_4 = io_tag_4; // @[S8DP1.scala 33:14:@665.4]
  assign mux_io_tag_5 = io_tag_5; // @[S8DP1.scala 33:14:@666.4]
  assign mux_io_tag_6 = io_tag_6; // @[S8DP1.scala 33:14:@667.4]
  assign mux_io_tag_7 = io_tag_7; // @[S8DP1.scala 33:14:@668.4]
  assign tag_change_clock = clock; // @[:@651.4]
  assign tag_change_reset = reset; // @[:@652.4]
  assign tag_change_io_tag_in_0 = io_tag_0; // @[S8DP1.scala 37:24:@674.4]
  assign tag_change_io_tag_in_1 = io_tag_1; // @[S8DP1.scala 37:24:@675.4]
  assign tag_change_io_tag_in_2 = io_tag_2; // @[S8DP1.scala 37:24:@676.4]
  assign tag_change_io_tag_in_3 = io_tag_3; // @[S8DP1.scala 37:24:@677.4]
  assign tag_change_io_tag_in_4 = io_tag_4; // @[S8DP1.scala 37:24:@678.4]
  assign tag_change_io_tag_in_5 = io_tag_5; // @[S8DP1.scala 37:24:@679.4]
  assign tag_change_io_tag_in_6 = io_tag_6; // @[S8DP1.scala 37:24:@680.4]
  assign tag_change_io_tag_in_7 = io_tag_7; // @[S8DP1.scala 37:24:@681.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  acc = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      acc <= 32'sh0;
    end else begin
      acc <= $signed(_GEN_1);
    end
  end
endmodule
module FF4( // @[:@7295.2]
  input clock, // @[:@7296.4]
  input reset, // @[:@7297.4]
  input [31:0] io_in_data_0_0, // @[:@7298.4]
  input [31:0] io_in_data_0_1, // @[:@7298.4]
  input [31:0] io_in_data_0_2, // @[:@7298.4]
  input [31:0] io_in_data_0_3, // @[:@7298.4]
  input [31:0] io_in_data_0_4, // @[:@7298.4]
  input [31:0] io_in_data_0_5, // @[:@7298.4]
  input [31:0] io_in_data_0_6, // @[:@7298.4]
  input [31:0] io_in_data_0_7, // @[:@7298.4]
  input [31:0] io_in_data_1_0, // @[:@7298.4]
  input [31:0] io_in_data_1_1, // @[:@7298.4]
  input [31:0] io_in_data_1_2, // @[:@7298.4]
  input [31:0] io_in_data_1_3, // @[:@7298.4]
  input [31:0] io_in_data_1_4, // @[:@7298.4]
  input [31:0] io_in_data_1_5, // @[:@7298.4]
  input [31:0] io_in_data_1_6, // @[:@7298.4]
  input [31:0] io_in_data_1_7, // @[:@7298.4]
  input [31:0] io_in_data_2_0, // @[:@7298.4]
  input [31:0] io_in_data_2_1, // @[:@7298.4]
  input [31:0] io_in_data_2_2, // @[:@7298.4]
  input [31:0] io_in_data_2_3, // @[:@7298.4]
  input [31:0] io_in_data_2_4, // @[:@7298.4]
  input [31:0] io_in_data_2_5, // @[:@7298.4]
  input [31:0] io_in_data_2_6, // @[:@7298.4]
  input [31:0] io_in_data_2_7, // @[:@7298.4]
  input [31:0] io_in_data_3_0, // @[:@7298.4]
  input [31:0] io_in_data_3_1, // @[:@7298.4]
  input [31:0] io_in_data_3_2, // @[:@7298.4]
  input [31:0] io_in_data_3_3, // @[:@7298.4]
  input [31:0] io_in_data_3_4, // @[:@7298.4]
  input [31:0] io_in_data_3_5, // @[:@7298.4]
  input [31:0] io_in_data_3_6, // @[:@7298.4]
  input [31:0] io_in_data_3_7, // @[:@7298.4]
  input io_in_tag_0_0, // @[:@7298.4]
  input io_in_tag_0_1, // @[:@7298.4]
  input io_in_tag_0_2, // @[:@7298.4]
  input io_in_tag_0_3, // @[:@7298.4]
  input io_in_tag_0_4, // @[:@7298.4]
  input io_in_tag_0_5, // @[:@7298.4]
  input io_in_tag_0_6, // @[:@7298.4]
  input io_in_tag_0_7, // @[:@7298.4]
  input io_in_tag_1_0, // @[:@7298.4]
  input io_in_tag_1_1, // @[:@7298.4]
  input io_in_tag_1_2, // @[:@7298.4]
  input io_in_tag_1_3, // @[:@7298.4]
  input io_in_tag_1_4, // @[:@7298.4]
  input io_in_tag_1_5, // @[:@7298.4]
  input io_in_tag_1_6, // @[:@7298.4]
  input io_in_tag_1_7, // @[:@7298.4]
  input io_in_tag_2_0, // @[:@7298.4]
  input io_in_tag_2_1, // @[:@7298.4]
  input io_in_tag_2_2, // @[:@7298.4]
  input io_in_tag_2_3, // @[:@7298.4]
  input io_in_tag_2_4, // @[:@7298.4]
  input io_in_tag_2_5, // @[:@7298.4]
  input io_in_tag_2_6, // @[:@7298.4]
  input io_in_tag_2_7, // @[:@7298.4]
  input io_in_tag_3_0, // @[:@7298.4]
  input io_in_tag_3_1, // @[:@7298.4]
  input io_in_tag_3_2, // @[:@7298.4]
  input io_in_tag_3_3, // @[:@7298.4]
  input io_in_tag_3_4, // @[:@7298.4]
  input io_in_tag_3_5, // @[:@7298.4]
  input io_in_tag_3_6, // @[:@7298.4]
  input io_in_tag_3_7, // @[:@7298.4]
  output [31:0] io_out_data_0_0, // @[:@7298.4]
  output [31:0] io_out_data_0_1, // @[:@7298.4]
  output [31:0] io_out_data_0_2, // @[:@7298.4]
  output [31:0] io_out_data_0_3, // @[:@7298.4]
  output [31:0] io_out_data_0_4, // @[:@7298.4]
  output [31:0] io_out_data_0_5, // @[:@7298.4]
  output [31:0] io_out_data_0_6, // @[:@7298.4]
  output [31:0] io_out_data_0_7, // @[:@7298.4]
  output [31:0] io_out_data_1_0, // @[:@7298.4]
  output [31:0] io_out_data_1_1, // @[:@7298.4]
  output [31:0] io_out_data_1_2, // @[:@7298.4]
  output [31:0] io_out_data_1_3, // @[:@7298.4]
  output [31:0] io_out_data_1_4, // @[:@7298.4]
  output [31:0] io_out_data_1_5, // @[:@7298.4]
  output [31:0] io_out_data_1_6, // @[:@7298.4]
  output [31:0] io_out_data_1_7, // @[:@7298.4]
  output [31:0] io_out_data_2_0, // @[:@7298.4]
  output [31:0] io_out_data_2_1, // @[:@7298.4]
  output [31:0] io_out_data_2_2, // @[:@7298.4]
  output [31:0] io_out_data_2_3, // @[:@7298.4]
  output [31:0] io_out_data_2_4, // @[:@7298.4]
  output [31:0] io_out_data_2_5, // @[:@7298.4]
  output [31:0] io_out_data_2_6, // @[:@7298.4]
  output [31:0] io_out_data_2_7, // @[:@7298.4]
  output [31:0] io_out_data_3_0, // @[:@7298.4]
  output [31:0] io_out_data_3_1, // @[:@7298.4]
  output [31:0] io_out_data_3_2, // @[:@7298.4]
  output [31:0] io_out_data_3_3, // @[:@7298.4]
  output [31:0] io_out_data_3_4, // @[:@7298.4]
  output [31:0] io_out_data_3_5, // @[:@7298.4]
  output [31:0] io_out_data_3_6, // @[:@7298.4]
  output [31:0] io_out_data_3_7, // @[:@7298.4]
  output io_out_tag_0_0, // @[:@7298.4]
  output io_out_tag_0_1, // @[:@7298.4]
  output io_out_tag_0_2, // @[:@7298.4]
  output io_out_tag_0_3, // @[:@7298.4]
  output io_out_tag_0_4, // @[:@7298.4]
  output io_out_tag_0_5, // @[:@7298.4]
  output io_out_tag_0_6, // @[:@7298.4]
  output io_out_tag_0_7, // @[:@7298.4]
  output io_out_tag_1_0, // @[:@7298.4]
  output io_out_tag_1_1, // @[:@7298.4]
  output io_out_tag_1_2, // @[:@7298.4]
  output io_out_tag_1_3, // @[:@7298.4]
  output io_out_tag_1_4, // @[:@7298.4]
  output io_out_tag_1_5, // @[:@7298.4]
  output io_out_tag_1_6, // @[:@7298.4]
  output io_out_tag_1_7, // @[:@7298.4]
  output io_out_tag_2_0, // @[:@7298.4]
  output io_out_tag_2_1, // @[:@7298.4]
  output io_out_tag_2_2, // @[:@7298.4]
  output io_out_tag_2_3, // @[:@7298.4]
  output io_out_tag_2_4, // @[:@7298.4]
  output io_out_tag_2_5, // @[:@7298.4]
  output io_out_tag_2_6, // @[:@7298.4]
  output io_out_tag_2_7, // @[:@7298.4]
  output io_out_tag_3_0, // @[:@7298.4]
  output io_out_tag_3_1, // @[:@7298.4]
  output io_out_tag_3_2, // @[:@7298.4]
  output io_out_tag_3_3, // @[:@7298.4]
  output io_out_tag_3_4, // @[:@7298.4]
  output io_out_tag_3_5, // @[:@7298.4]
  output io_out_tag_3_6, // @[:@7298.4]
  output io_out_tag_3_7 // @[:@7298.4]
);
  reg [31:0] data_0_0; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_0;
  reg [31:0] data_0_1; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_1;
  reg [31:0] data_0_2; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_2;
  reg [31:0] data_0_3; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_3;
  reg [31:0] data_0_4; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_4;
  reg [31:0] data_0_5; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_5;
  reg [31:0] data_0_6; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_6;
  reg [31:0] data_0_7; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_7;
  reg [31:0] data_1_0; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_8;
  reg [31:0] data_1_1; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_9;
  reg [31:0] data_1_2; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_10;
  reg [31:0] data_1_3; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_11;
  reg [31:0] data_1_4; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_12;
  reg [31:0] data_1_5; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_13;
  reg [31:0] data_1_6; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_14;
  reg [31:0] data_1_7; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_15;
  reg [31:0] data_2_0; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_16;
  reg [31:0] data_2_1; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_17;
  reg [31:0] data_2_2; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_18;
  reg [31:0] data_2_3; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_19;
  reg [31:0] data_2_4; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_20;
  reg [31:0] data_2_5; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_21;
  reg [31:0] data_2_6; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_22;
  reg [31:0] data_2_7; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_23;
  reg [31:0] data_3_0; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_24;
  reg [31:0] data_3_1; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_25;
  reg [31:0] data_3_2; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_26;
  reg [31:0] data_3_3; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_27;
  reg [31:0] data_3_4; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_28;
  reg [31:0] data_3_5; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_29;
  reg [31:0] data_3_6; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_30;
  reg [31:0] data_3_7; // @[FF4.scala 63:21:@7369.4]
  reg [31:0] _RAND_31;
  reg tag_0_0; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_32;
  reg tag_0_1; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_33;
  reg tag_0_2; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_34;
  reg tag_0_3; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_35;
  reg tag_0_4; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_36;
  reg tag_0_5; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_37;
  reg tag_0_6; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_38;
  reg tag_0_7; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_39;
  reg tag_1_0; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_40;
  reg tag_1_1; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_41;
  reg tag_1_2; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_42;
  reg tag_1_3; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_43;
  reg tag_1_4; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_44;
  reg tag_1_5; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_45;
  reg tag_1_6; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_46;
  reg tag_1_7; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_47;
  reg tag_2_0; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_48;
  reg tag_2_1; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_49;
  reg tag_2_2; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_50;
  reg tag_2_3; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_51;
  reg tag_2_4; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_52;
  reg tag_2_5; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_53;
  reg tag_2_6; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_54;
  reg tag_2_7; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_55;
  reg tag_3_0; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_56;
  reg tag_3_1; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_57;
  reg tag_3_2; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_58;
  reg tag_3_3; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_59;
  reg tag_3_4; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_60;
  reg tag_3_5; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_61;
  reg tag_3_6; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_62;
  reg tag_3_7; // @[FF4.scala 64:20:@7439.4]
  reg [31:0] _RAND_63;
  assign io_out_data_0_0 = data_0_0; // @[FF4.scala 69:15:@7504.4]
  assign io_out_data_0_1 = data_0_1; // @[FF4.scala 69:15:@7505.4]
  assign io_out_data_0_2 = data_0_2; // @[FF4.scala 69:15:@7506.4]
  assign io_out_data_0_3 = data_0_3; // @[FF4.scala 69:15:@7507.4]
  assign io_out_data_0_4 = data_0_4; // @[FF4.scala 69:15:@7508.4]
  assign io_out_data_0_5 = data_0_5; // @[FF4.scala 69:15:@7509.4]
  assign io_out_data_0_6 = data_0_6; // @[FF4.scala 69:15:@7510.4]
  assign io_out_data_0_7 = data_0_7; // @[FF4.scala 69:15:@7511.4]
  assign io_out_data_1_0 = data_1_0; // @[FF4.scala 69:15:@7512.4]
  assign io_out_data_1_1 = data_1_1; // @[FF4.scala 69:15:@7513.4]
  assign io_out_data_1_2 = data_1_2; // @[FF4.scala 69:15:@7514.4]
  assign io_out_data_1_3 = data_1_3; // @[FF4.scala 69:15:@7515.4]
  assign io_out_data_1_4 = data_1_4; // @[FF4.scala 69:15:@7516.4]
  assign io_out_data_1_5 = data_1_5; // @[FF4.scala 69:15:@7517.4]
  assign io_out_data_1_6 = data_1_6; // @[FF4.scala 69:15:@7518.4]
  assign io_out_data_1_7 = data_1_7; // @[FF4.scala 69:15:@7519.4]
  assign io_out_data_2_0 = data_2_0; // @[FF4.scala 69:15:@7520.4]
  assign io_out_data_2_1 = data_2_1; // @[FF4.scala 69:15:@7521.4]
  assign io_out_data_2_2 = data_2_2; // @[FF4.scala 69:15:@7522.4]
  assign io_out_data_2_3 = data_2_3; // @[FF4.scala 69:15:@7523.4]
  assign io_out_data_2_4 = data_2_4; // @[FF4.scala 69:15:@7524.4]
  assign io_out_data_2_5 = data_2_5; // @[FF4.scala 69:15:@7525.4]
  assign io_out_data_2_6 = data_2_6; // @[FF4.scala 69:15:@7526.4]
  assign io_out_data_2_7 = data_2_7; // @[FF4.scala 69:15:@7527.4]
  assign io_out_data_3_0 = data_3_0; // @[FF4.scala 69:15:@7528.4]
  assign io_out_data_3_1 = data_3_1; // @[FF4.scala 69:15:@7529.4]
  assign io_out_data_3_2 = data_3_2; // @[FF4.scala 69:15:@7530.4]
  assign io_out_data_3_3 = data_3_3; // @[FF4.scala 69:15:@7531.4]
  assign io_out_data_3_4 = data_3_4; // @[FF4.scala 69:15:@7532.4]
  assign io_out_data_3_5 = data_3_5; // @[FF4.scala 69:15:@7533.4]
  assign io_out_data_3_6 = data_3_6; // @[FF4.scala 69:15:@7534.4]
  assign io_out_data_3_7 = data_3_7; // @[FF4.scala 69:15:@7535.4]
  assign io_out_tag_0_0 = tag_0_0; // @[FF4.scala 70:14:@7536.4]
  assign io_out_tag_0_1 = tag_0_1; // @[FF4.scala 70:14:@7537.4]
  assign io_out_tag_0_2 = tag_0_2; // @[FF4.scala 70:14:@7538.4]
  assign io_out_tag_0_3 = tag_0_3; // @[FF4.scala 70:14:@7539.4]
  assign io_out_tag_0_4 = tag_0_4; // @[FF4.scala 70:14:@7540.4]
  assign io_out_tag_0_5 = tag_0_5; // @[FF4.scala 70:14:@7541.4]
  assign io_out_tag_0_6 = tag_0_6; // @[FF4.scala 70:14:@7542.4]
  assign io_out_tag_0_7 = tag_0_7; // @[FF4.scala 70:14:@7543.4]
  assign io_out_tag_1_0 = tag_1_0; // @[FF4.scala 70:14:@7544.4]
  assign io_out_tag_1_1 = tag_1_1; // @[FF4.scala 70:14:@7545.4]
  assign io_out_tag_1_2 = tag_1_2; // @[FF4.scala 70:14:@7546.4]
  assign io_out_tag_1_3 = tag_1_3; // @[FF4.scala 70:14:@7547.4]
  assign io_out_tag_1_4 = tag_1_4; // @[FF4.scala 70:14:@7548.4]
  assign io_out_tag_1_5 = tag_1_5; // @[FF4.scala 70:14:@7549.4]
  assign io_out_tag_1_6 = tag_1_6; // @[FF4.scala 70:14:@7550.4]
  assign io_out_tag_1_7 = tag_1_7; // @[FF4.scala 70:14:@7551.4]
  assign io_out_tag_2_0 = tag_2_0; // @[FF4.scala 70:14:@7552.4]
  assign io_out_tag_2_1 = tag_2_1; // @[FF4.scala 70:14:@7553.4]
  assign io_out_tag_2_2 = tag_2_2; // @[FF4.scala 70:14:@7554.4]
  assign io_out_tag_2_3 = tag_2_3; // @[FF4.scala 70:14:@7555.4]
  assign io_out_tag_2_4 = tag_2_4; // @[FF4.scala 70:14:@7556.4]
  assign io_out_tag_2_5 = tag_2_5; // @[FF4.scala 70:14:@7557.4]
  assign io_out_tag_2_6 = tag_2_6; // @[FF4.scala 70:14:@7558.4]
  assign io_out_tag_2_7 = tag_2_7; // @[FF4.scala 70:14:@7559.4]
  assign io_out_tag_3_0 = tag_3_0; // @[FF4.scala 70:14:@7560.4]
  assign io_out_tag_3_1 = tag_3_1; // @[FF4.scala 70:14:@7561.4]
  assign io_out_tag_3_2 = tag_3_2; // @[FF4.scala 70:14:@7562.4]
  assign io_out_tag_3_3 = tag_3_3; // @[FF4.scala 70:14:@7563.4]
  assign io_out_tag_3_4 = tag_3_4; // @[FF4.scala 70:14:@7564.4]
  assign io_out_tag_3_5 = tag_3_5; // @[FF4.scala 70:14:@7565.4]
  assign io_out_tag_3_6 = tag_3_6; // @[FF4.scala 70:14:@7566.4]
  assign io_out_tag_3_7 = tag_3_7; // @[FF4.scala 70:14:@7567.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  data_0_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  data_0_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  data_0_2 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  data_0_3 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  data_0_4 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  data_0_5 = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  data_0_6 = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  data_0_7 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  data_1_0 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  data_1_1 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  data_1_2 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  data_1_3 = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  data_1_4 = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  data_1_5 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  data_1_6 = _RAND_14[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  data_1_7 = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  data_2_0 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  data_2_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  data_2_2 = _RAND_18[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  data_2_3 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  data_2_4 = _RAND_20[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  data_2_5 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  data_2_6 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  data_2_7 = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  data_3_0 = _RAND_24[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  data_3_1 = _RAND_25[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  data_3_2 = _RAND_26[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  data_3_3 = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  data_3_4 = _RAND_28[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  data_3_5 = _RAND_29[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  data_3_6 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  data_3_7 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_32 = {1{$random}};
  tag_0_0 = _RAND_32[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_33 = {1{$random}};
  tag_0_1 = _RAND_33[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_34 = {1{$random}};
  tag_0_2 = _RAND_34[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_35 = {1{$random}};
  tag_0_3 = _RAND_35[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_36 = {1{$random}};
  tag_0_4 = _RAND_36[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_37 = {1{$random}};
  tag_0_5 = _RAND_37[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_38 = {1{$random}};
  tag_0_6 = _RAND_38[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_39 = {1{$random}};
  tag_0_7 = _RAND_39[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_40 = {1{$random}};
  tag_1_0 = _RAND_40[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_41 = {1{$random}};
  tag_1_1 = _RAND_41[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_42 = {1{$random}};
  tag_1_2 = _RAND_42[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_43 = {1{$random}};
  tag_1_3 = _RAND_43[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_44 = {1{$random}};
  tag_1_4 = _RAND_44[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_45 = {1{$random}};
  tag_1_5 = _RAND_45[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_46 = {1{$random}};
  tag_1_6 = _RAND_46[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_47 = {1{$random}};
  tag_1_7 = _RAND_47[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_48 = {1{$random}};
  tag_2_0 = _RAND_48[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_49 = {1{$random}};
  tag_2_1 = _RAND_49[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_50 = {1{$random}};
  tag_2_2 = _RAND_50[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_51 = {1{$random}};
  tag_2_3 = _RAND_51[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_52 = {1{$random}};
  tag_2_4 = _RAND_52[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_53 = {1{$random}};
  tag_2_5 = _RAND_53[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_54 = {1{$random}};
  tag_2_6 = _RAND_54[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_55 = {1{$random}};
  tag_2_7 = _RAND_55[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_56 = {1{$random}};
  tag_3_0 = _RAND_56[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_57 = {1{$random}};
  tag_3_1 = _RAND_57[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_58 = {1{$random}};
  tag_3_2 = _RAND_58[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_59 = {1{$random}};
  tag_3_3 = _RAND_59[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_60 = {1{$random}};
  tag_3_4 = _RAND_60[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_61 = {1{$random}};
  tag_3_5 = _RAND_61[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_62 = {1{$random}};
  tag_3_6 = _RAND_62[0:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_63 = {1{$random}};
  tag_3_7 = _RAND_63[0:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      data_0_0 <= 32'sh0;
    end else begin
      data_0_0 <= io_in_data_0_0;
    end
    if (reset) begin
      data_0_1 <= 32'sh0;
    end else begin
      data_0_1 <= io_in_data_0_1;
    end
    if (reset) begin
      data_0_2 <= 32'sh0;
    end else begin
      data_0_2 <= io_in_data_0_2;
    end
    if (reset) begin
      data_0_3 <= 32'sh0;
    end else begin
      data_0_3 <= io_in_data_0_3;
    end
    if (reset) begin
      data_0_4 <= 32'sh0;
    end else begin
      data_0_4 <= io_in_data_0_4;
    end
    if (reset) begin
      data_0_5 <= 32'sh0;
    end else begin
      data_0_5 <= io_in_data_0_5;
    end
    if (reset) begin
      data_0_6 <= 32'sh0;
    end else begin
      data_0_6 <= io_in_data_0_6;
    end
    if (reset) begin
      data_0_7 <= 32'sh0;
    end else begin
      data_0_7 <= io_in_data_0_7;
    end
    if (reset) begin
      data_1_0 <= 32'sh0;
    end else begin
      data_1_0 <= io_in_data_1_0;
    end
    if (reset) begin
      data_1_1 <= 32'sh0;
    end else begin
      data_1_1 <= io_in_data_1_1;
    end
    if (reset) begin
      data_1_2 <= 32'sh0;
    end else begin
      data_1_2 <= io_in_data_1_2;
    end
    if (reset) begin
      data_1_3 <= 32'sh0;
    end else begin
      data_1_3 <= io_in_data_1_3;
    end
    if (reset) begin
      data_1_4 <= 32'sh0;
    end else begin
      data_1_4 <= io_in_data_1_4;
    end
    if (reset) begin
      data_1_5 <= 32'sh0;
    end else begin
      data_1_5 <= io_in_data_1_5;
    end
    if (reset) begin
      data_1_6 <= 32'sh0;
    end else begin
      data_1_6 <= io_in_data_1_6;
    end
    if (reset) begin
      data_1_7 <= 32'sh0;
    end else begin
      data_1_7 <= io_in_data_1_7;
    end
    if (reset) begin
      data_2_0 <= 32'sh0;
    end else begin
      data_2_0 <= io_in_data_2_0;
    end
    if (reset) begin
      data_2_1 <= 32'sh0;
    end else begin
      data_2_1 <= io_in_data_2_1;
    end
    if (reset) begin
      data_2_2 <= 32'sh0;
    end else begin
      data_2_2 <= io_in_data_2_2;
    end
    if (reset) begin
      data_2_3 <= 32'sh0;
    end else begin
      data_2_3 <= io_in_data_2_3;
    end
    if (reset) begin
      data_2_4 <= 32'sh0;
    end else begin
      data_2_4 <= io_in_data_2_4;
    end
    if (reset) begin
      data_2_5 <= 32'sh0;
    end else begin
      data_2_5 <= io_in_data_2_5;
    end
    if (reset) begin
      data_2_6 <= 32'sh0;
    end else begin
      data_2_6 <= io_in_data_2_6;
    end
    if (reset) begin
      data_2_7 <= 32'sh0;
    end else begin
      data_2_7 <= io_in_data_2_7;
    end
    if (reset) begin
      data_3_0 <= 32'sh0;
    end else begin
      data_3_0 <= io_in_data_3_0;
    end
    if (reset) begin
      data_3_1 <= 32'sh0;
    end else begin
      data_3_1 <= io_in_data_3_1;
    end
    if (reset) begin
      data_3_2 <= 32'sh0;
    end else begin
      data_3_2 <= io_in_data_3_2;
    end
    if (reset) begin
      data_3_3 <= 32'sh0;
    end else begin
      data_3_3 <= io_in_data_3_3;
    end
    if (reset) begin
      data_3_4 <= 32'sh0;
    end else begin
      data_3_4 <= io_in_data_3_4;
    end
    if (reset) begin
      data_3_5 <= 32'sh0;
    end else begin
      data_3_5 <= io_in_data_3_5;
    end
    if (reset) begin
      data_3_6 <= 32'sh0;
    end else begin
      data_3_6 <= io_in_data_3_6;
    end
    if (reset) begin
      data_3_7 <= 32'sh0;
    end else begin
      data_3_7 <= io_in_data_3_7;
    end
    if (reset) begin
      tag_0_0 <= 1'h0;
    end else begin
      tag_0_0 <= io_in_tag_0_0;
    end
    if (reset) begin
      tag_0_1 <= 1'h0;
    end else begin
      tag_0_1 <= io_in_tag_0_1;
    end
    if (reset) begin
      tag_0_2 <= 1'h0;
    end else begin
      tag_0_2 <= io_in_tag_0_2;
    end
    if (reset) begin
      tag_0_3 <= 1'h0;
    end else begin
      tag_0_3 <= io_in_tag_0_3;
    end
    if (reset) begin
      tag_0_4 <= 1'h0;
    end else begin
      tag_0_4 <= io_in_tag_0_4;
    end
    if (reset) begin
      tag_0_5 <= 1'h0;
    end else begin
      tag_0_5 <= io_in_tag_0_5;
    end
    if (reset) begin
      tag_0_6 <= 1'h0;
    end else begin
      tag_0_6 <= io_in_tag_0_6;
    end
    if (reset) begin
      tag_0_7 <= 1'h0;
    end else begin
      tag_0_7 <= io_in_tag_0_7;
    end
    if (reset) begin
      tag_1_0 <= 1'h0;
    end else begin
      tag_1_0 <= io_in_tag_1_0;
    end
    if (reset) begin
      tag_1_1 <= 1'h0;
    end else begin
      tag_1_1 <= io_in_tag_1_1;
    end
    if (reset) begin
      tag_1_2 <= 1'h0;
    end else begin
      tag_1_2 <= io_in_tag_1_2;
    end
    if (reset) begin
      tag_1_3 <= 1'h0;
    end else begin
      tag_1_3 <= io_in_tag_1_3;
    end
    if (reset) begin
      tag_1_4 <= 1'h0;
    end else begin
      tag_1_4 <= io_in_tag_1_4;
    end
    if (reset) begin
      tag_1_5 <= 1'h0;
    end else begin
      tag_1_5 <= io_in_tag_1_5;
    end
    if (reset) begin
      tag_1_6 <= 1'h0;
    end else begin
      tag_1_6 <= io_in_tag_1_6;
    end
    if (reset) begin
      tag_1_7 <= 1'h0;
    end else begin
      tag_1_7 <= io_in_tag_1_7;
    end
    if (reset) begin
      tag_2_0 <= 1'h0;
    end else begin
      tag_2_0 <= io_in_tag_2_0;
    end
    if (reset) begin
      tag_2_1 <= 1'h0;
    end else begin
      tag_2_1 <= io_in_tag_2_1;
    end
    if (reset) begin
      tag_2_2 <= 1'h0;
    end else begin
      tag_2_2 <= io_in_tag_2_2;
    end
    if (reset) begin
      tag_2_3 <= 1'h0;
    end else begin
      tag_2_3 <= io_in_tag_2_3;
    end
    if (reset) begin
      tag_2_4 <= 1'h0;
    end else begin
      tag_2_4 <= io_in_tag_2_4;
    end
    if (reset) begin
      tag_2_5 <= 1'h0;
    end else begin
      tag_2_5 <= io_in_tag_2_5;
    end
    if (reset) begin
      tag_2_6 <= 1'h0;
    end else begin
      tag_2_6 <= io_in_tag_2_6;
    end
    if (reset) begin
      tag_2_7 <= 1'h0;
    end else begin
      tag_2_7 <= io_in_tag_2_7;
    end
    if (reset) begin
      tag_3_0 <= 1'h0;
    end else begin
      tag_3_0 <= io_in_tag_3_0;
    end
    if (reset) begin
      tag_3_1 <= 1'h0;
    end else begin
      tag_3_1 <= io_in_tag_3_1;
    end
    if (reset) begin
      tag_3_2 <= 1'h0;
    end else begin
      tag_3_2 <= io_in_tag_3_2;
    end
    if (reset) begin
      tag_3_3 <= 1'h0;
    end else begin
      tag_3_3 <= io_in_tag_3_3;
    end
    if (reset) begin
      tag_3_4 <= 1'h0;
    end else begin
      tag_3_4 <= io_in_tag_3_4;
    end
    if (reset) begin
      tag_3_5 <= 1'h0;
    end else begin
      tag_3_5 <= io_in_tag_3_5;
    end
    if (reset) begin
      tag_3_6 <= 1'h0;
    end else begin
      tag_3_6 <= io_in_tag_3_6;
    end
    if (reset) begin
      tag_3_7 <= 1'h0;
    end else begin
      tag_3_7 <= io_in_tag_3_7;
    end
  end
endmodule
module FF8( // @[:@7843.2]
  input clock, // @[:@7844.4]
  input reset, // @[:@7845.4]
  input [31:0] io_in_data_0_0, // @[:@7846.4]
  input [31:0] io_in_data_0_1, // @[:@7846.4]
  input [31:0] io_in_data_0_2, // @[:@7846.4]
  input [31:0] io_in_data_0_3, // @[:@7846.4]
  input [31:0] io_in_data_0_4, // @[:@7846.4]
  input [31:0] io_in_data_0_5, // @[:@7846.4]
  input [31:0] io_in_data_0_6, // @[:@7846.4]
  input [31:0] io_in_data_0_7, // @[:@7846.4]
  input [31:0] io_in_data_1_0, // @[:@7846.4]
  input [31:0] io_in_data_1_1, // @[:@7846.4]
  input [31:0] io_in_data_1_2, // @[:@7846.4]
  input [31:0] io_in_data_1_3, // @[:@7846.4]
  input [31:0] io_in_data_1_4, // @[:@7846.4]
  input [31:0] io_in_data_1_5, // @[:@7846.4]
  input [31:0] io_in_data_1_6, // @[:@7846.4]
  input [31:0] io_in_data_1_7, // @[:@7846.4]
  output [31:0] io_out_data_0_0, // @[:@7846.4]
  output [31:0] io_out_data_0_1, // @[:@7846.4]
  output [31:0] io_out_data_0_2, // @[:@7846.4]
  output [31:0] io_out_data_0_3, // @[:@7846.4]
  output [31:0] io_out_data_0_4, // @[:@7846.4]
  output [31:0] io_out_data_0_5, // @[:@7846.4]
  output [31:0] io_out_data_0_6, // @[:@7846.4]
  output [31:0] io_out_data_0_7, // @[:@7846.4]
  output [31:0] io_out_data_1_0, // @[:@7846.4]
  output [31:0] io_out_data_1_1, // @[:@7846.4]
  output [31:0] io_out_data_1_2, // @[:@7846.4]
  output [31:0] io_out_data_1_3, // @[:@7846.4]
  output [31:0] io_out_data_1_4, // @[:@7846.4]
  output [31:0] io_out_data_1_5, // @[:@7846.4]
  output [31:0] io_out_data_1_6, // @[:@7846.4]
  output [31:0] io_out_data_1_7 // @[:@7846.4]
);
  reg [31:0] data_0_0; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_0;
  reg [31:0] data_0_1; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_1;
  reg [31:0] data_0_2; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_2;
  reg [31:0] data_0_3; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_3;
  reg [31:0] data_0_4; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_4;
  reg [31:0] data_0_5; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_5;
  reg [31:0] data_0_6; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_6;
  reg [31:0] data_0_7; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_7;
  reg [31:0] data_1_0; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_8;
  reg [31:0] data_1_1; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_9;
  reg [31:0] data_1_2; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_10;
  reg [31:0] data_1_3; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_11;
  reg [31:0] data_1_4; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_12;
  reg [31:0] data_1_5; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_13;
  reg [31:0] data_1_6; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_14;
  reg [31:0] data_1_7; // @[FF8.scala 72:21:@7883.4]
  reg [31:0] _RAND_15;
  assign io_out_data_0_0 = data_0_0; // @[FF8.scala 74:15:@7900.4]
  assign io_out_data_0_1 = data_0_1; // @[FF8.scala 74:15:@7901.4]
  assign io_out_data_0_2 = data_0_2; // @[FF8.scala 74:15:@7902.4]
  assign io_out_data_0_3 = data_0_3; // @[FF8.scala 74:15:@7903.4]
  assign io_out_data_0_4 = data_0_4; // @[FF8.scala 74:15:@7904.4]
  assign io_out_data_0_5 = data_0_5; // @[FF8.scala 74:15:@7905.4]
  assign io_out_data_0_6 = data_0_6; // @[FF8.scala 74:15:@7906.4]
  assign io_out_data_0_7 = data_0_7; // @[FF8.scala 74:15:@7907.4]
  assign io_out_data_1_0 = data_1_0; // @[FF8.scala 74:15:@7908.4]
  assign io_out_data_1_1 = data_1_1; // @[FF8.scala 74:15:@7909.4]
  assign io_out_data_1_2 = data_1_2; // @[FF8.scala 74:15:@7910.4]
  assign io_out_data_1_3 = data_1_3; // @[FF8.scala 74:15:@7911.4]
  assign io_out_data_1_4 = data_1_4; // @[FF8.scala 74:15:@7912.4]
  assign io_out_data_1_5 = data_1_5; // @[FF8.scala 74:15:@7913.4]
  assign io_out_data_1_6 = data_1_6; // @[FF8.scala 74:15:@7914.4]
  assign io_out_data_1_7 = data_1_7; // @[FF8.scala 74:15:@7915.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  data_0_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  data_0_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  data_0_2 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  data_0_3 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  data_0_4 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  data_0_5 = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  data_0_6 = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  data_0_7 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  data_1_0 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  data_1_1 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  data_1_2 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  data_1_3 = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  data_1_4 = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  data_1_5 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  data_1_6 = _RAND_14[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  data_1_7 = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      data_0_0 <= 32'sh0;
    end else begin
      data_0_0 <= io_in_data_0_0;
    end
    if (reset) begin
      data_0_1 <= 32'sh0;
    end else begin
      data_0_1 <= io_in_data_0_1;
    end
    if (reset) begin
      data_0_2 <= 32'sh0;
    end else begin
      data_0_2 <= io_in_data_0_2;
    end
    if (reset) begin
      data_0_3 <= 32'sh0;
    end else begin
      data_0_3 <= io_in_data_0_3;
    end
    if (reset) begin
      data_0_4 <= 32'sh0;
    end else begin
      data_0_4 <= io_in_data_0_4;
    end
    if (reset) begin
      data_0_5 <= 32'sh0;
    end else begin
      data_0_5 <= io_in_data_0_5;
    end
    if (reset) begin
      data_0_6 <= 32'sh0;
    end else begin
      data_0_6 <= io_in_data_0_6;
    end
    if (reset) begin
      data_0_7 <= 32'sh0;
    end else begin
      data_0_7 <= io_in_data_0_7;
    end
    if (reset) begin
      data_1_0 <= 32'sh0;
    end else begin
      data_1_0 <= io_in_data_1_0;
    end
    if (reset) begin
      data_1_1 <= 32'sh0;
    end else begin
      data_1_1 <= io_in_data_1_1;
    end
    if (reset) begin
      data_1_2 <= 32'sh0;
    end else begin
      data_1_2 <= io_in_data_1_2;
    end
    if (reset) begin
      data_1_3 <= 32'sh0;
    end else begin
      data_1_3 <= io_in_data_1_3;
    end
    if (reset) begin
      data_1_4 <= 32'sh0;
    end else begin
      data_1_4 <= io_in_data_1_4;
    end
    if (reset) begin
      data_1_5 <= 32'sh0;
    end else begin
      data_1_5 <= io_in_data_1_5;
    end
    if (reset) begin
      data_1_6 <= 32'sh0;
    end else begin
      data_1_6 <= io_in_data_1_6;
    end
    if (reset) begin
      data_1_7 <= 32'sh0;
    end else begin
      data_1_7 <= io_in_data_1_7;
    end
  end
endmodule
module STA_VDBB( // @[:@8687.2]
  input clock, // @[:@8688.4]
  input reset, // @[:@8689.4]
  input [31:0] io_in_A_0_0, // @[:@8690.4]
  input [31:0] io_in_A_0_1, // @[:@8690.4]
  input [31:0] io_in_A_0_2, // @[:@8690.4]
  input [31:0] io_in_A_0_3, // @[:@8690.4]
  input [31:0] io_in_A_0_4, // @[:@8690.4]
  input [31:0] io_in_A_0_5, // @[:@8690.4]
  input [31:0] io_in_A_0_6, // @[:@8690.4]
  input [31:0] io_in_A_0_7, // @[:@8690.4]
  input [31:0] io_in_A_0_8, // @[:@8690.4]
  input [31:0] io_in_A_0_9, // @[:@8690.4]
  input [31:0] io_in_A_0_10, // @[:@8690.4]
  input [31:0] io_in_A_0_11, // @[:@8690.4]
  input [31:0] io_in_A_0_12, // @[:@8690.4]
  input [31:0] io_in_A_0_13, // @[:@8690.4]
  input [31:0] io_in_A_0_14, // @[:@8690.4]
  input [31:0] io_in_A_0_15, // @[:@8690.4]
  input [31:0] io_in_A_1_0, // @[:@8690.4]
  input [31:0] io_in_A_1_1, // @[:@8690.4]
  input [31:0] io_in_A_1_2, // @[:@8690.4]
  input [31:0] io_in_A_1_3, // @[:@8690.4]
  input [31:0] io_in_A_1_4, // @[:@8690.4]
  input [31:0] io_in_A_1_5, // @[:@8690.4]
  input [31:0] io_in_A_1_6, // @[:@8690.4]
  input [31:0] io_in_A_1_7, // @[:@8690.4]
  input [31:0] io_in_A_1_8, // @[:@8690.4]
  input [31:0] io_in_A_1_9, // @[:@8690.4]
  input [31:0] io_in_A_1_10, // @[:@8690.4]
  input [31:0] io_in_A_1_11, // @[:@8690.4]
  input [31:0] io_in_A_1_12, // @[:@8690.4]
  input [31:0] io_in_A_1_13, // @[:@8690.4]
  input [31:0] io_in_A_1_14, // @[:@8690.4]
  input [31:0] io_in_A_1_15, // @[:@8690.4]
  input [31:0] io_in_A_2_0, // @[:@8690.4]
  input [31:0] io_in_A_2_1, // @[:@8690.4]
  input [31:0] io_in_A_2_2, // @[:@8690.4]
  input [31:0] io_in_A_2_3, // @[:@8690.4]
  input [31:0] io_in_A_2_4, // @[:@8690.4]
  input [31:0] io_in_A_2_5, // @[:@8690.4]
  input [31:0] io_in_A_2_6, // @[:@8690.4]
  input [31:0] io_in_A_2_7, // @[:@8690.4]
  input [31:0] io_in_A_2_8, // @[:@8690.4]
  input [31:0] io_in_A_2_9, // @[:@8690.4]
  input [31:0] io_in_A_2_10, // @[:@8690.4]
  input [31:0] io_in_A_2_11, // @[:@8690.4]
  input [31:0] io_in_A_2_12, // @[:@8690.4]
  input [31:0] io_in_A_2_13, // @[:@8690.4]
  input [31:0] io_in_A_2_14, // @[:@8690.4]
  input [31:0] io_in_A_2_15, // @[:@8690.4]
  input [31:0] io_in_A_3_0, // @[:@8690.4]
  input [31:0] io_in_A_3_1, // @[:@8690.4]
  input [31:0] io_in_A_3_2, // @[:@8690.4]
  input [31:0] io_in_A_3_3, // @[:@8690.4]
  input [31:0] io_in_A_3_4, // @[:@8690.4]
  input [31:0] io_in_A_3_5, // @[:@8690.4]
  input [31:0] io_in_A_3_6, // @[:@8690.4]
  input [31:0] io_in_A_3_7, // @[:@8690.4]
  input [31:0] io_in_A_3_8, // @[:@8690.4]
  input [31:0] io_in_A_3_9, // @[:@8690.4]
  input [31:0] io_in_A_3_10, // @[:@8690.4]
  input [31:0] io_in_A_3_11, // @[:@8690.4]
  input [31:0] io_in_A_3_12, // @[:@8690.4]
  input [31:0] io_in_A_3_13, // @[:@8690.4]
  input [31:0] io_in_A_3_14, // @[:@8690.4]
  input [31:0] io_in_A_3_15, // @[:@8690.4]
  input [31:0] io_in_B_0_0, // @[:@8690.4]
  input [31:0] io_in_B_0_1, // @[:@8690.4]
  input [31:0] io_in_B_0_2, // @[:@8690.4]
  input [31:0] io_in_B_0_3, // @[:@8690.4]
  input [31:0] io_in_B_0_4, // @[:@8690.4]
  input [31:0] io_in_B_0_5, // @[:@8690.4]
  input [31:0] io_in_B_0_6, // @[:@8690.4]
  input [31:0] io_in_B_0_7, // @[:@8690.4]
  input [31:0] io_in_B_0_8, // @[:@8690.4]
  input [31:0] io_in_B_0_9, // @[:@8690.4]
  input [31:0] io_in_B_0_10, // @[:@8690.4]
  input [31:0] io_in_B_0_11, // @[:@8690.4]
  input [31:0] io_in_B_0_12, // @[:@8690.4]
  input [31:0] io_in_B_0_13, // @[:@8690.4]
  input [31:0] io_in_B_0_14, // @[:@8690.4]
  input [31:0] io_in_B_0_15, // @[:@8690.4]
  input [31:0] io_in_B_1_0, // @[:@8690.4]
  input [31:0] io_in_B_1_1, // @[:@8690.4]
  input [31:0] io_in_B_1_2, // @[:@8690.4]
  input [31:0] io_in_B_1_3, // @[:@8690.4]
  input [31:0] io_in_B_1_4, // @[:@8690.4]
  input [31:0] io_in_B_1_5, // @[:@8690.4]
  input [31:0] io_in_B_1_6, // @[:@8690.4]
  input [31:0] io_in_B_1_7, // @[:@8690.4]
  input [31:0] io_in_B_1_8, // @[:@8690.4]
  input [31:0] io_in_B_1_9, // @[:@8690.4]
  input [31:0] io_in_B_1_10, // @[:@8690.4]
  input [31:0] io_in_B_1_11, // @[:@8690.4]
  input [31:0] io_in_B_1_12, // @[:@8690.4]
  input [31:0] io_in_B_1_13, // @[:@8690.4]
  input [31:0] io_in_B_1_14, // @[:@8690.4]
  input [31:0] io_in_B_1_15, // @[:@8690.4]
  input [31:0] io_in_B_2_0, // @[:@8690.4]
  input [31:0] io_in_B_2_1, // @[:@8690.4]
  input [31:0] io_in_B_2_2, // @[:@8690.4]
  input [31:0] io_in_B_2_3, // @[:@8690.4]
  input [31:0] io_in_B_2_4, // @[:@8690.4]
  input [31:0] io_in_B_2_5, // @[:@8690.4]
  input [31:0] io_in_B_2_6, // @[:@8690.4]
  input [31:0] io_in_B_2_7, // @[:@8690.4]
  input [31:0] io_in_B_2_8, // @[:@8690.4]
  input [31:0] io_in_B_2_9, // @[:@8690.4]
  input [31:0] io_in_B_2_10, // @[:@8690.4]
  input [31:0] io_in_B_2_11, // @[:@8690.4]
  input [31:0] io_in_B_2_12, // @[:@8690.4]
  input [31:0] io_in_B_2_13, // @[:@8690.4]
  input [31:0] io_in_B_2_14, // @[:@8690.4]
  input [31:0] io_in_B_2_15, // @[:@8690.4]
  input [31:0] io_in_B_3_0, // @[:@8690.4]
  input [31:0] io_in_B_3_1, // @[:@8690.4]
  input [31:0] io_in_B_3_2, // @[:@8690.4]
  input [31:0] io_in_B_3_3, // @[:@8690.4]
  input [31:0] io_in_B_3_4, // @[:@8690.4]
  input [31:0] io_in_B_3_5, // @[:@8690.4]
  input [31:0] io_in_B_3_6, // @[:@8690.4]
  input [31:0] io_in_B_3_7, // @[:@8690.4]
  input [31:0] io_in_B_3_8, // @[:@8690.4]
  input [31:0] io_in_B_3_9, // @[:@8690.4]
  input [31:0] io_in_B_3_10, // @[:@8690.4]
  input [31:0] io_in_B_3_11, // @[:@8690.4]
  input [31:0] io_in_B_3_12, // @[:@8690.4]
  input [31:0] io_in_B_3_13, // @[:@8690.4]
  input [31:0] io_in_B_3_14, // @[:@8690.4]
  input [31:0] io_in_B_3_15, // @[:@8690.4]
  input [31:0] io_in_B_4_0, // @[:@8690.4]
  input [31:0] io_in_B_4_1, // @[:@8690.4]
  input [31:0] io_in_B_4_2, // @[:@8690.4]
  input [31:0] io_in_B_4_3, // @[:@8690.4]
  input [31:0] io_in_B_4_4, // @[:@8690.4]
  input [31:0] io_in_B_4_5, // @[:@8690.4]
  input [31:0] io_in_B_4_6, // @[:@8690.4]
  input [31:0] io_in_B_4_7, // @[:@8690.4]
  input [31:0] io_in_B_4_8, // @[:@8690.4]
  input [31:0] io_in_B_4_9, // @[:@8690.4]
  input [31:0] io_in_B_4_10, // @[:@8690.4]
  input [31:0] io_in_B_4_11, // @[:@8690.4]
  input [31:0] io_in_B_4_12, // @[:@8690.4]
  input [31:0] io_in_B_4_13, // @[:@8690.4]
  input [31:0] io_in_B_4_14, // @[:@8690.4]
  input [31:0] io_in_B_4_15, // @[:@8690.4]
  input [31:0] io_in_B_5_0, // @[:@8690.4]
  input [31:0] io_in_B_5_1, // @[:@8690.4]
  input [31:0] io_in_B_5_2, // @[:@8690.4]
  input [31:0] io_in_B_5_3, // @[:@8690.4]
  input [31:0] io_in_B_5_4, // @[:@8690.4]
  input [31:0] io_in_B_5_5, // @[:@8690.4]
  input [31:0] io_in_B_5_6, // @[:@8690.4]
  input [31:0] io_in_B_5_7, // @[:@8690.4]
  input [31:0] io_in_B_5_8, // @[:@8690.4]
  input [31:0] io_in_B_5_9, // @[:@8690.4]
  input [31:0] io_in_B_5_10, // @[:@8690.4]
  input [31:0] io_in_B_5_11, // @[:@8690.4]
  input [31:0] io_in_B_5_12, // @[:@8690.4]
  input [31:0] io_in_B_5_13, // @[:@8690.4]
  input [31:0] io_in_B_5_14, // @[:@8690.4]
  input [31:0] io_in_B_5_15, // @[:@8690.4]
  input [31:0] io_in_B_6_0, // @[:@8690.4]
  input [31:0] io_in_B_6_1, // @[:@8690.4]
  input [31:0] io_in_B_6_2, // @[:@8690.4]
  input [31:0] io_in_B_6_3, // @[:@8690.4]
  input [31:0] io_in_B_6_4, // @[:@8690.4]
  input [31:0] io_in_B_6_5, // @[:@8690.4]
  input [31:0] io_in_B_6_6, // @[:@8690.4]
  input [31:0] io_in_B_6_7, // @[:@8690.4]
  input [31:0] io_in_B_6_8, // @[:@8690.4]
  input [31:0] io_in_B_6_9, // @[:@8690.4]
  input [31:0] io_in_B_6_10, // @[:@8690.4]
  input [31:0] io_in_B_6_11, // @[:@8690.4]
  input [31:0] io_in_B_6_12, // @[:@8690.4]
  input [31:0] io_in_B_6_13, // @[:@8690.4]
  input [31:0] io_in_B_6_14, // @[:@8690.4]
  input [31:0] io_in_B_6_15, // @[:@8690.4]
  input [31:0] io_in_B_7_0, // @[:@8690.4]
  input [31:0] io_in_B_7_1, // @[:@8690.4]
  input [31:0] io_in_B_7_2, // @[:@8690.4]
  input [31:0] io_in_B_7_3, // @[:@8690.4]
  input [31:0] io_in_B_7_4, // @[:@8690.4]
  input [31:0] io_in_B_7_5, // @[:@8690.4]
  input [31:0] io_in_B_7_6, // @[:@8690.4]
  input [31:0] io_in_B_7_7, // @[:@8690.4]
  input [31:0] io_in_B_7_8, // @[:@8690.4]
  input [31:0] io_in_B_7_9, // @[:@8690.4]
  input [31:0] io_in_B_7_10, // @[:@8690.4]
  input [31:0] io_in_B_7_11, // @[:@8690.4]
  input [31:0] io_in_B_7_12, // @[:@8690.4]
  input [31:0] io_in_B_7_13, // @[:@8690.4]
  input [31:0] io_in_B_7_14, // @[:@8690.4]
  input [31:0] io_in_B_7_15, // @[:@8690.4]
  output [31:0] io_out_C_0_0, // @[:@8690.4]
  output [31:0] io_out_C_0_1, // @[:@8690.4]
  output [31:0] io_out_C_0_2, // @[:@8690.4]
  output [31:0] io_out_C_0_3, // @[:@8690.4]
  output [31:0] io_out_C_0_4, // @[:@8690.4]
  output [31:0] io_out_C_0_5, // @[:@8690.4]
  output [31:0] io_out_C_0_6, // @[:@8690.4]
  output [31:0] io_out_C_0_7, // @[:@8690.4]
  output [31:0] io_out_C_1_0, // @[:@8690.4]
  output [31:0] io_out_C_1_1, // @[:@8690.4]
  output [31:0] io_out_C_1_2, // @[:@8690.4]
  output [31:0] io_out_C_1_3, // @[:@8690.4]
  output [31:0] io_out_C_1_4, // @[:@8690.4]
  output [31:0] io_out_C_1_5, // @[:@8690.4]
  output [31:0] io_out_C_1_6, // @[:@8690.4]
  output [31:0] io_out_C_1_7, // @[:@8690.4]
  output [31:0] io_out_C_2_0, // @[:@8690.4]
  output [31:0] io_out_C_2_1, // @[:@8690.4]
  output [31:0] io_out_C_2_2, // @[:@8690.4]
  output [31:0] io_out_C_2_3, // @[:@8690.4]
  output [31:0] io_out_C_2_4, // @[:@8690.4]
  output [31:0] io_out_C_2_5, // @[:@8690.4]
  output [31:0] io_out_C_2_6, // @[:@8690.4]
  output [31:0] io_out_C_2_7, // @[:@8690.4]
  output [31:0] io_out_C_3_0, // @[:@8690.4]
  output [31:0] io_out_C_3_1, // @[:@8690.4]
  output [31:0] io_out_C_3_2, // @[:@8690.4]
  output [31:0] io_out_C_3_3, // @[:@8690.4]
  output [31:0] io_out_C_3_4, // @[:@8690.4]
  output [31:0] io_out_C_3_5, // @[:@8690.4]
  output [31:0] io_out_C_3_6, // @[:@8690.4]
  output [31:0] io_out_C_3_7 // @[:@8690.4]
);
  wire tag_clock; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_reset; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_0; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_1; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_2; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_3; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_4; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_5; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_io_out_tag_6; // @[STA_VDBB.scala 51:39:@8692.4]
  wire tag_1_clock; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_reset; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_0; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_1; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_2; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_3; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_4; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_5; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_1_io_out_tag_6; // @[STA_VDBB.scala 51:39:@8695.4]
  wire tag_2_clock; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_reset; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_0; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_1; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_2; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_3; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_4; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_5; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_2_io_out_tag_6; // @[STA_VDBB.scala 51:39:@8698.4]
  wire tag_3_clock; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_reset; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_0; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_1; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_2; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_3; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_4; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_5; // @[STA_VDBB.scala 51:39:@8701.4]
  wire tag_3_io_out_tag_6; // @[STA_VDBB.scala 51:39:@8701.4]
  wire [31:0] MUX8_io_int_in_0; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_1; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_2; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_3; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_4; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_5; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_6; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_int_in_7; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_0; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_1; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_2; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_3; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_4; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_5; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_6; // @[STA_VDBB.scala 52:36:@8773.4]
  wire MUX8_io_tag_7; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_io_choice; // @[STA_VDBB.scala 52:36:@8773.4]
  wire [31:0] MUX8_1_io_int_in_0; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_1; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_2; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_3; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_4; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_5; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_6; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_int_in_7; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_0; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_1; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_2; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_3; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_4; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_5; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_6; // @[STA_VDBB.scala 52:36:@8776.4]
  wire MUX8_1_io_tag_7; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_1_io_choice; // @[STA_VDBB.scala 52:36:@8776.4]
  wire [31:0] MUX8_2_io_int_in_0; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_1; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_2; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_3; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_4; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_5; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_6; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_int_in_7; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_0; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_1; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_2; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_3; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_4; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_5; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_6; // @[STA_VDBB.scala 52:36:@8779.4]
  wire MUX8_2_io_tag_7; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_2_io_choice; // @[STA_VDBB.scala 52:36:@8779.4]
  wire [31:0] MUX8_3_io_int_in_0; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_1; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_2; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_3; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_4; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_5; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_6; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_int_in_7; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_0; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_1; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_2; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_3; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_4; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_5; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_6; // @[STA_VDBB.scala 52:36:@8782.4]
  wire MUX8_3_io_tag_7; // @[STA_VDBB.scala 52:36:@8782.4]
  wire [31:0] MUX8_3_io_choice; // @[STA_VDBB.scala 52:36:@8782.4]
  wire S8DP1_clock; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_reset; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_int_in_B; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_0; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_1; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_2; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_3; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_4; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_5; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_6; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_tag_7; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8854.4]
  wire [31:0] S8DP1_io_result; // @[STA_VDBB.scala 55:44:@8854.4]
  wire S8DP1_1_clock; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_reset; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_int_in_B; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_0; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_1; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_2; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_3; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_4; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_5; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_6; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_tag_7; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_1_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8857.4]
  wire [31:0] S8DP1_1_io_result; // @[STA_VDBB.scala 55:44:@8857.4]
  wire S8DP1_2_clock; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_reset; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_int_in_B; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_0; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_1; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_2; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_3; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_4; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_5; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_6; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_tag_7; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_2_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8860.4]
  wire [31:0] S8DP1_2_io_result; // @[STA_VDBB.scala 55:44:@8860.4]
  wire S8DP1_3_clock; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_reset; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_int_in_B; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_0; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_1; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_2; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_3; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_4; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_5; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_6; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_tag_7; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_3_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8863.4]
  wire [31:0] S8DP1_3_io_result; // @[STA_VDBB.scala 55:44:@8863.4]
  wire S8DP1_4_clock; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_reset; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_int_in_B; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_0; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_1; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_2; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_3; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_4; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_5; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_6; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_tag_7; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_4_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8866.4]
  wire [31:0] S8DP1_4_io_result; // @[STA_VDBB.scala 55:44:@8866.4]
  wire S8DP1_5_clock; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_reset; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_int_in_B; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_0; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_1; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_2; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_3; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_4; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_5; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_6; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_tag_7; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_5_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8869.4]
  wire [31:0] S8DP1_5_io_result; // @[STA_VDBB.scala 55:44:@8869.4]
  wire S8DP1_6_clock; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_reset; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_int_in_B; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_0; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_1; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_2; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_3; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_4; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_5; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_6; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_tag_7; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_6_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8872.4]
  wire [31:0] S8DP1_6_io_result; // @[STA_VDBB.scala 55:44:@8872.4]
  wire S8DP1_7_clock; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_reset; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_0; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_1; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_2; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_3; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_4; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_5; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_6; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_A_7; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_int_in_B; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_0; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_1; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_2; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_3; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_4; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_5; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_6; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_tag_7; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_0; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_1; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_2; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_3; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_4; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_5; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_6; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_7_io_out_tag_7; // @[STA_VDBB.scala 55:44:@8875.4]
  wire [31:0] S8DP1_7_io_result; // @[STA_VDBB.scala 55:44:@8875.4]
  wire S8DP1_8_clock; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_reset; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_int_in_B; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_0; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_1; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_2; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_3; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_4; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_5; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_6; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_tag_7; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_8_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9087.4]
  wire [31:0] S8DP1_8_io_result; // @[STA_VDBB.scala 56:44:@9087.4]
  wire S8DP1_9_clock; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_reset; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_int_in_B; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_0; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_1; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_2; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_3; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_4; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_5; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_6; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_tag_7; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_9_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9090.4]
  wire [31:0] S8DP1_9_io_result; // @[STA_VDBB.scala 56:44:@9090.4]
  wire S8DP1_10_clock; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_reset; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_int_in_B; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_0; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_1; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_2; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_3; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_4; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_5; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_6; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_tag_7; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_10_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9093.4]
  wire [31:0] S8DP1_10_io_result; // @[STA_VDBB.scala 56:44:@9093.4]
  wire S8DP1_11_clock; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_reset; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_int_in_B; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_0; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_1; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_2; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_3; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_4; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_5; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_6; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_tag_7; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_11_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9096.4]
  wire [31:0] S8DP1_11_io_result; // @[STA_VDBB.scala 56:44:@9096.4]
  wire S8DP1_12_clock; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_reset; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_int_in_B; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_0; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_1; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_2; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_3; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_4; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_5; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_6; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_tag_7; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_12_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9099.4]
  wire [31:0] S8DP1_12_io_result; // @[STA_VDBB.scala 56:44:@9099.4]
  wire S8DP1_13_clock; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_reset; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_int_in_B; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_0; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_1; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_2; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_3; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_4; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_5; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_6; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_tag_7; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_13_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9102.4]
  wire [31:0] S8DP1_13_io_result; // @[STA_VDBB.scala 56:44:@9102.4]
  wire S8DP1_14_clock; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_reset; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_int_in_B; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_0; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_1; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_2; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_3; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_4; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_5; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_6; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_tag_7; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_14_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9105.4]
  wire [31:0] S8DP1_14_io_result; // @[STA_VDBB.scala 56:44:@9105.4]
  wire S8DP1_15_clock; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_reset; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_0; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_1; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_2; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_3; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_4; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_5; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_6; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_A_7; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_int_in_B; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_0; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_1; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_2; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_3; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_4; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_5; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_6; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_tag_7; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_0; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_1; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_2; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_3; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_4; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_5; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_6; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_15_io_out_tag_7; // @[STA_VDBB.scala 56:44:@9108.4]
  wire [31:0] S8DP1_15_io_result; // @[STA_VDBB.scala 56:44:@9108.4]
  wire S8DP1_16_clock; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_reset; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_int_in_B; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_0; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_1; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_2; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_3; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_4; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_5; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_6; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_tag_7; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_16_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9320.4]
  wire [31:0] S8DP1_16_io_result; // @[STA_VDBB.scala 57:44:@9320.4]
  wire S8DP1_17_clock; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_reset; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_int_in_B; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_0; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_1; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_2; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_3; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_4; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_5; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_6; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_tag_7; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_17_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9323.4]
  wire [31:0] S8DP1_17_io_result; // @[STA_VDBB.scala 57:44:@9323.4]
  wire S8DP1_18_clock; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_reset; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_int_in_B; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_0; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_1; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_2; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_3; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_4; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_5; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_6; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_tag_7; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_18_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9326.4]
  wire [31:0] S8DP1_18_io_result; // @[STA_VDBB.scala 57:44:@9326.4]
  wire S8DP1_19_clock; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_reset; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_int_in_B; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_0; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_1; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_2; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_3; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_4; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_5; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_6; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_tag_7; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_19_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9329.4]
  wire [31:0] S8DP1_19_io_result; // @[STA_VDBB.scala 57:44:@9329.4]
  wire S8DP1_20_clock; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_reset; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_int_in_B; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_0; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_1; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_2; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_3; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_4; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_5; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_6; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_tag_7; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_20_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9332.4]
  wire [31:0] S8DP1_20_io_result; // @[STA_VDBB.scala 57:44:@9332.4]
  wire S8DP1_21_clock; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_reset; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_int_in_B; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_0; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_1; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_2; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_3; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_4; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_5; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_6; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_tag_7; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_21_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9335.4]
  wire [31:0] S8DP1_21_io_result; // @[STA_VDBB.scala 57:44:@9335.4]
  wire S8DP1_22_clock; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_reset; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_int_in_B; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_0; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_1; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_2; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_3; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_4; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_5; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_6; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_tag_7; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_22_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9338.4]
  wire [31:0] S8DP1_22_io_result; // @[STA_VDBB.scala 57:44:@9338.4]
  wire S8DP1_23_clock; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_reset; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_0; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_1; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_2; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_3; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_4; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_5; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_6; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_A_7; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_int_in_B; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_0; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_1; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_2; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_3; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_4; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_5; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_6; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_tag_7; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_0; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_1; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_2; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_3; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_4; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_5; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_6; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_23_io_out_tag_7; // @[STA_VDBB.scala 57:44:@9341.4]
  wire [31:0] S8DP1_23_io_result; // @[STA_VDBB.scala 57:44:@9341.4]
  wire S8DP1_24_clock; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_reset; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_int_in_B; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_0; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_1; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_2; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_3; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_4; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_5; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_6; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_tag_7; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_24_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9553.4]
  wire [31:0] S8DP1_24_io_result; // @[STA_VDBB.scala 58:44:@9553.4]
  wire S8DP1_25_clock; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_reset; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_int_in_B; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_0; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_1; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_2; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_3; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_4; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_5; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_6; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_tag_7; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_25_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9556.4]
  wire [31:0] S8DP1_25_io_result; // @[STA_VDBB.scala 58:44:@9556.4]
  wire S8DP1_26_clock; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_reset; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_int_in_B; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_0; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_1; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_2; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_3; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_4; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_5; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_6; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_tag_7; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_26_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9559.4]
  wire [31:0] S8DP1_26_io_result; // @[STA_VDBB.scala 58:44:@9559.4]
  wire S8DP1_27_clock; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_reset; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_int_in_B; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_0; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_1; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_2; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_3; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_4; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_5; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_6; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_tag_7; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_27_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9562.4]
  wire [31:0] S8DP1_27_io_result; // @[STA_VDBB.scala 58:44:@9562.4]
  wire S8DP1_28_clock; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_reset; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_int_in_B; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_0; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_1; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_2; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_3; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_4; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_5; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_6; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_tag_7; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_28_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9565.4]
  wire [31:0] S8DP1_28_io_result; // @[STA_VDBB.scala 58:44:@9565.4]
  wire S8DP1_29_clock; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_reset; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_int_in_B; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_0; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_1; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_2; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_3; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_4; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_5; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_6; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_tag_7; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_29_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9568.4]
  wire [31:0] S8DP1_29_io_result; // @[STA_VDBB.scala 58:44:@9568.4]
  wire S8DP1_30_clock; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_reset; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_int_in_B; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_0; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_1; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_2; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_3; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_4; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_5; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_6; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_tag_7; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_30_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9571.4]
  wire [31:0] S8DP1_30_io_result; // @[STA_VDBB.scala 58:44:@9571.4]
  wire S8DP1_31_clock; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_reset; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_0; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_1; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_2; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_3; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_4; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_5; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_6; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_A_7; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_int_in_B; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_0; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_1; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_2; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_3; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_4; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_5; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_6; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_tag_7; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_0; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_1; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_2; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_3; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_4; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_5; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_6; // @[STA_VDBB.scala 58:44:@9574.4]
  wire S8DP1_31_io_out_tag_7; // @[STA_VDBB.scala 58:44:@9574.4]
  wire [31:0] S8DP1_31_io_result; // @[STA_VDBB.scala 58:44:@9574.4]
  wire ffb1_clock; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_reset; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_0_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_1_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_2_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_in_data_3_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_0_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_1_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_2_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_in_tag_3_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_0_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_1_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_2_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire [31:0] ffb1_io_out_data_3_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_0_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_1_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_2_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_0; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_1; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_2; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_3; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_4; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_5; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_6; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb1_io_out_tag_3_7; // @[STA_VDBB.scala 68:20:@9786.4]
  wire ffb2_clock; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_reset; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_0_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_1_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_2_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_in_data_3_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_0_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_1_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_2_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_in_tag_3_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_0_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_1_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_2_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire [31:0] ffb2_io_out_data_3_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_0_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_1_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_2_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_0; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_1; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_2; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_3; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_4; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_5; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_6; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffb2_io_out_tag_3_7; // @[STA_VDBB.scala 69:20:@9789.4]
  wire ffa1_clock; // @[STA_VDBB.scala 71:20:@9792.4]
  wire ffa1_reset; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_0; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_1; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_2; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_3; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_4; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_5; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_6; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_0_7; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_0; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_1; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_2; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_3; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_4; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_5; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_6; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_in_data_1_7; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_0; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_1; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_2; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_3; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_4; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_5; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_6; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_0_7; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_0; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_1; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_2; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_3; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_4; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_5; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_6; // @[STA_VDBB.scala 71:20:@9792.4]
  wire [31:0] ffa1_io_out_data_1_7; // @[STA_VDBB.scala 71:20:@9792.4]
  wire ff00_clock; // @[STA_VDBB.scala 72:20:@9795.4]
  wire ff00_reset; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_0; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_1; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_2; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_3; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_4; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_5; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_6; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_0_7; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_0; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_1; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_2; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_3; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_4; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_5; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_6; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_in_data_1_7; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_0; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_1; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_2; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_3; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_4; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_5; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_6; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_0_7; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_0; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_1; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_2; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_3; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_4; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_5; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_6; // @[STA_VDBB.scala 72:20:@9795.4]
  wire [31:0] ff00_io_out_data_1_7; // @[STA_VDBB.scala 72:20:@9795.4]
  wire ff01_clock; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_reset; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_0_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_1_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_2_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_in_data_3_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_0_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_1_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_2_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_in_tag_3_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_0_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_1_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_2_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire [31:0] ff01_io_out_data_3_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_0_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_1_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_2_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_0; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_1; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_2; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_3; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_4; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_5; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_6; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff01_io_out_tag_3_7; // @[STA_VDBB.scala 74:20:@9798.4]
  wire ff10_clock; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_reset; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_0_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_1_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_2_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_in_data_3_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_0_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_1_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_2_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_in_tag_3_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_0_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_1_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_2_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire [31:0] ff10_io_out_data_3_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_0_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_1_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_2_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_0; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_1; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_2; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_3; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_4; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_5; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_6; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ff10_io_out_tag_3_7; // @[STA_VDBB.scala 75:20:@9801.4]
  wire ffa2_clock; // @[STA_VDBB.scala 77:20:@9804.4]
  wire ffa2_reset; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_0; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_1; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_2; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_3; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_4; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_5; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_6; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_0_7; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_0; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_1; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_2; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_3; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_4; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_5; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_6; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_in_data_1_7; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_0; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_1; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_2; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_3; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_4; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_5; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_6; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_0_7; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_0; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_1; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_2; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_3; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_4; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_5; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_6; // @[STA_VDBB.scala 77:20:@9804.4]
  wire [31:0] ffa2_io_out_data_1_7; // @[STA_VDBB.scala 77:20:@9804.4]
  wire ff11_clock; // @[STA_VDBB.scala 78:20:@9807.4]
  wire ff11_reset; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_0; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_1; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_2; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_3; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_4; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_5; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_6; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_0_7; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_0; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_1; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_2; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_3; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_4; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_5; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_6; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_in_data_1_7; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_0; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_1; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_2; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_3; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_4; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_5; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_6; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_0_7; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_0; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_1; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_2; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_3; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_4; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_5; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_6; // @[STA_VDBB.scala 78:20:@9807.4]
  wire [31:0] ff11_io_out_data_1_7; // @[STA_VDBB.scala 78:20:@9807.4]
  reg [31:0] out_result_0_0; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_0;
  reg [31:0] out_result_0_1; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_1;
  reg [31:0] out_result_0_2; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_2;
  reg [31:0] out_result_0_3; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_3;
  reg [31:0] out_result_0_4; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_4;
  reg [31:0] out_result_0_5; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_5;
  reg [31:0] out_result_0_6; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_6;
  reg [31:0] out_result_0_7; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_7;
  reg [31:0] out_result_1_0; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_8;
  reg [31:0] out_result_1_1; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_9;
  reg [31:0] out_result_1_2; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_10;
  reg [31:0] out_result_1_3; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_11;
  reg [31:0] out_result_1_4; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_12;
  reg [31:0] out_result_1_5; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_13;
  reg [31:0] out_result_1_6; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_14;
  reg [31:0] out_result_1_7; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_15;
  reg [31:0] out_result_2_0; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_16;
  reg [31:0] out_result_2_1; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_17;
  reg [31:0] out_result_2_2; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_18;
  reg [31:0] out_result_2_3; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_19;
  reg [31:0] out_result_2_4; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_20;
  reg [31:0] out_result_2_5; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_21;
  reg [31:0] out_result_2_6; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_22;
  reg [31:0] out_result_2_7; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_23;
  reg [31:0] out_result_3_0; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_24;
  reg [31:0] out_result_3_1; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_25;
  reg [31:0] out_result_3_2; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_26;
  reg [31:0] out_result_3_3; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_27;
  reg [31:0] out_result_3_4; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_28;
  reg [31:0] out_result_3_5; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_29;
  reg [31:0] out_result_3_6; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_30;
  reg [31:0] out_result_3_7; // @[STA_VDBB.scala 346:27:@27809.4]
  reg [31:0] _RAND_31;
  wire [31:0] S8DP1s_0_0_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8879.4]
  wire [31:0] S8DP1s_0_1_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8905.4]
  wire [31:0] S8DP1s_0_2_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8931.4]
  wire [31:0] S8DP1s_0_3_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8957.4]
  wire [31:0] S8DP1s_0_4_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8983.4]
  wire [31:0] S8DP1s_0_5_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9009.4]
  wire [31:0] S8DP1s_0_6_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9035.4]
  wire [31:0] S8DP1s_0_7_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9061.4]
  wire [31:0] S8DP1s_1_0_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9112.4]
  wire [31:0] S8DP1s_1_1_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9138.4]
  wire [31:0] S8DP1s_1_2_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9164.4]
  wire [31:0] S8DP1s_1_3_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9190.4]
  wire [31:0] S8DP1s_1_4_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9216.4]
  wire [31:0] S8DP1s_1_5_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9242.4]
  wire [31:0] S8DP1s_1_6_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9268.4]
  wire [31:0] S8DP1s_1_7_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9294.4]
  wire [31:0] S8DP1s_2_0_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9345.4]
  wire [31:0] S8DP1s_2_1_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9371.4]
  wire [31:0] S8DP1s_2_2_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9397.4]
  wire [31:0] S8DP1s_2_3_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9423.4]
  wire [31:0] S8DP1s_2_4_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9449.4]
  wire [31:0] S8DP1s_2_5_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9475.4]
  wire [31:0] S8DP1s_2_6_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9501.4]
  wire [31:0] S8DP1s_2_7_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9527.4]
  wire [31:0] S8DP1s_3_0_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9578.4]
  wire [31:0] S8DP1s_3_1_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9604.4]
  wire [31:0] S8DP1s_3_2_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9630.4]
  wire [31:0] S8DP1s_3_3_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9656.4]
  wire [31:0] S8DP1s_3_4_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9682.4]
  wire [31:0] S8DP1s_3_5_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9708.4]
  wire [31:0] S8DP1s_3_6_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9734.4]
  wire [31:0] S8DP1s_3_7_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9760.4]
  tag tag( // @[STA_VDBB.scala 51:39:@8692.4]
    .clock(tag_clock),
    .reset(tag_reset),
    .io_out_tag_0(tag_io_out_tag_0),
    .io_out_tag_1(tag_io_out_tag_1),
    .io_out_tag_2(tag_io_out_tag_2),
    .io_out_tag_3(tag_io_out_tag_3),
    .io_out_tag_4(tag_io_out_tag_4),
    .io_out_tag_5(tag_io_out_tag_5),
    .io_out_tag_6(tag_io_out_tag_6)
  );
  tag tag_1( // @[STA_VDBB.scala 51:39:@8695.4]
    .clock(tag_1_clock),
    .reset(tag_1_reset),
    .io_out_tag_0(tag_1_io_out_tag_0),
    .io_out_tag_1(tag_1_io_out_tag_1),
    .io_out_tag_2(tag_1_io_out_tag_2),
    .io_out_tag_3(tag_1_io_out_tag_3),
    .io_out_tag_4(tag_1_io_out_tag_4),
    .io_out_tag_5(tag_1_io_out_tag_5),
    .io_out_tag_6(tag_1_io_out_tag_6)
  );
  tag tag_2( // @[STA_VDBB.scala 51:39:@8698.4]
    .clock(tag_2_clock),
    .reset(tag_2_reset),
    .io_out_tag_0(tag_2_io_out_tag_0),
    .io_out_tag_1(tag_2_io_out_tag_1),
    .io_out_tag_2(tag_2_io_out_tag_2),
    .io_out_tag_3(tag_2_io_out_tag_3),
    .io_out_tag_4(tag_2_io_out_tag_4),
    .io_out_tag_5(tag_2_io_out_tag_5),
    .io_out_tag_6(tag_2_io_out_tag_6)
  );
  tag tag_3( // @[STA_VDBB.scala 51:39:@8701.4]
    .clock(tag_3_clock),
    .reset(tag_3_reset),
    .io_out_tag_0(tag_3_io_out_tag_0),
    .io_out_tag_1(tag_3_io_out_tag_1),
    .io_out_tag_2(tag_3_io_out_tag_2),
    .io_out_tag_3(tag_3_io_out_tag_3),
    .io_out_tag_4(tag_3_io_out_tag_4),
    .io_out_tag_5(tag_3_io_out_tag_5),
    .io_out_tag_6(tag_3_io_out_tag_6)
  );
  MUX8 MUX8( // @[STA_VDBB.scala 52:36:@8773.4]
    .io_int_in_0(MUX8_io_int_in_0),
    .io_int_in_1(MUX8_io_int_in_1),
    .io_int_in_2(MUX8_io_int_in_2),
    .io_int_in_3(MUX8_io_int_in_3),
    .io_int_in_4(MUX8_io_int_in_4),
    .io_int_in_5(MUX8_io_int_in_5),
    .io_int_in_6(MUX8_io_int_in_6),
    .io_int_in_7(MUX8_io_int_in_7),
    .io_tag_0(MUX8_io_tag_0),
    .io_tag_1(MUX8_io_tag_1),
    .io_tag_2(MUX8_io_tag_2),
    .io_tag_3(MUX8_io_tag_3),
    .io_tag_4(MUX8_io_tag_4),
    .io_tag_5(MUX8_io_tag_5),
    .io_tag_6(MUX8_io_tag_6),
    .io_tag_7(MUX8_io_tag_7),
    .io_choice(MUX8_io_choice)
  );
  MUX8 MUX8_1( // @[STA_VDBB.scala 52:36:@8776.4]
    .io_int_in_0(MUX8_1_io_int_in_0),
    .io_int_in_1(MUX8_1_io_int_in_1),
    .io_int_in_2(MUX8_1_io_int_in_2),
    .io_int_in_3(MUX8_1_io_int_in_3),
    .io_int_in_4(MUX8_1_io_int_in_4),
    .io_int_in_5(MUX8_1_io_int_in_5),
    .io_int_in_6(MUX8_1_io_int_in_6),
    .io_int_in_7(MUX8_1_io_int_in_7),
    .io_tag_0(MUX8_1_io_tag_0),
    .io_tag_1(MUX8_1_io_tag_1),
    .io_tag_2(MUX8_1_io_tag_2),
    .io_tag_3(MUX8_1_io_tag_3),
    .io_tag_4(MUX8_1_io_tag_4),
    .io_tag_5(MUX8_1_io_tag_5),
    .io_tag_6(MUX8_1_io_tag_6),
    .io_tag_7(MUX8_1_io_tag_7),
    .io_choice(MUX8_1_io_choice)
  );
  MUX8 MUX8_2( // @[STA_VDBB.scala 52:36:@8779.4]
    .io_int_in_0(MUX8_2_io_int_in_0),
    .io_int_in_1(MUX8_2_io_int_in_1),
    .io_int_in_2(MUX8_2_io_int_in_2),
    .io_int_in_3(MUX8_2_io_int_in_3),
    .io_int_in_4(MUX8_2_io_int_in_4),
    .io_int_in_5(MUX8_2_io_int_in_5),
    .io_int_in_6(MUX8_2_io_int_in_6),
    .io_int_in_7(MUX8_2_io_int_in_7),
    .io_tag_0(MUX8_2_io_tag_0),
    .io_tag_1(MUX8_2_io_tag_1),
    .io_tag_2(MUX8_2_io_tag_2),
    .io_tag_3(MUX8_2_io_tag_3),
    .io_tag_4(MUX8_2_io_tag_4),
    .io_tag_5(MUX8_2_io_tag_5),
    .io_tag_6(MUX8_2_io_tag_6),
    .io_tag_7(MUX8_2_io_tag_7),
    .io_choice(MUX8_2_io_choice)
  );
  MUX8 MUX8_3( // @[STA_VDBB.scala 52:36:@8782.4]
    .io_int_in_0(MUX8_3_io_int_in_0),
    .io_int_in_1(MUX8_3_io_int_in_1),
    .io_int_in_2(MUX8_3_io_int_in_2),
    .io_int_in_3(MUX8_3_io_int_in_3),
    .io_int_in_4(MUX8_3_io_int_in_4),
    .io_int_in_5(MUX8_3_io_int_in_5),
    .io_int_in_6(MUX8_3_io_int_in_6),
    .io_int_in_7(MUX8_3_io_int_in_7),
    .io_tag_0(MUX8_3_io_tag_0),
    .io_tag_1(MUX8_3_io_tag_1),
    .io_tag_2(MUX8_3_io_tag_2),
    .io_tag_3(MUX8_3_io_tag_3),
    .io_tag_4(MUX8_3_io_tag_4),
    .io_tag_5(MUX8_3_io_tag_5),
    .io_tag_6(MUX8_3_io_tag_6),
    .io_tag_7(MUX8_3_io_tag_7),
    .io_choice(MUX8_3_io_choice)
  );
  S8DP1 S8DP1( // @[STA_VDBB.scala 55:44:@8854.4]
    .clock(S8DP1_clock),
    .reset(S8DP1_reset),
    .io_int_in_A_0(S8DP1_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_io_int_in_A_7),
    .io_int_in_B(S8DP1_io_int_in_B),
    .io_tag_0(S8DP1_io_tag_0),
    .io_tag_1(S8DP1_io_tag_1),
    .io_tag_2(S8DP1_io_tag_2),
    .io_tag_3(S8DP1_io_tag_3),
    .io_tag_4(S8DP1_io_tag_4),
    .io_tag_5(S8DP1_io_tag_5),
    .io_tag_6(S8DP1_io_tag_6),
    .io_tag_7(S8DP1_io_tag_7),
    .io_out_tag_0(S8DP1_io_out_tag_0),
    .io_out_tag_1(S8DP1_io_out_tag_1),
    .io_out_tag_2(S8DP1_io_out_tag_2),
    .io_out_tag_3(S8DP1_io_out_tag_3),
    .io_out_tag_4(S8DP1_io_out_tag_4),
    .io_out_tag_5(S8DP1_io_out_tag_5),
    .io_out_tag_6(S8DP1_io_out_tag_6),
    .io_out_tag_7(S8DP1_io_out_tag_7),
    .io_result(S8DP1_io_result)
  );
  S8DP1 S8DP1_1( // @[STA_VDBB.scala 55:44:@8857.4]
    .clock(S8DP1_1_clock),
    .reset(S8DP1_1_reset),
    .io_int_in_A_0(S8DP1_1_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_1_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_1_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_1_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_1_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_1_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_1_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_1_io_int_in_A_7),
    .io_int_in_B(S8DP1_1_io_int_in_B),
    .io_tag_0(S8DP1_1_io_tag_0),
    .io_tag_1(S8DP1_1_io_tag_1),
    .io_tag_2(S8DP1_1_io_tag_2),
    .io_tag_3(S8DP1_1_io_tag_3),
    .io_tag_4(S8DP1_1_io_tag_4),
    .io_tag_5(S8DP1_1_io_tag_5),
    .io_tag_6(S8DP1_1_io_tag_6),
    .io_tag_7(S8DP1_1_io_tag_7),
    .io_out_tag_0(S8DP1_1_io_out_tag_0),
    .io_out_tag_1(S8DP1_1_io_out_tag_1),
    .io_out_tag_2(S8DP1_1_io_out_tag_2),
    .io_out_tag_3(S8DP1_1_io_out_tag_3),
    .io_out_tag_4(S8DP1_1_io_out_tag_4),
    .io_out_tag_5(S8DP1_1_io_out_tag_5),
    .io_out_tag_6(S8DP1_1_io_out_tag_6),
    .io_out_tag_7(S8DP1_1_io_out_tag_7),
    .io_result(S8DP1_1_io_result)
  );
  S8DP1 S8DP1_2( // @[STA_VDBB.scala 55:44:@8860.4]
    .clock(S8DP1_2_clock),
    .reset(S8DP1_2_reset),
    .io_int_in_A_0(S8DP1_2_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_2_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_2_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_2_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_2_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_2_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_2_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_2_io_int_in_A_7),
    .io_int_in_B(S8DP1_2_io_int_in_B),
    .io_tag_0(S8DP1_2_io_tag_0),
    .io_tag_1(S8DP1_2_io_tag_1),
    .io_tag_2(S8DP1_2_io_tag_2),
    .io_tag_3(S8DP1_2_io_tag_3),
    .io_tag_4(S8DP1_2_io_tag_4),
    .io_tag_5(S8DP1_2_io_tag_5),
    .io_tag_6(S8DP1_2_io_tag_6),
    .io_tag_7(S8DP1_2_io_tag_7),
    .io_out_tag_0(S8DP1_2_io_out_tag_0),
    .io_out_tag_1(S8DP1_2_io_out_tag_1),
    .io_out_tag_2(S8DP1_2_io_out_tag_2),
    .io_out_tag_3(S8DP1_2_io_out_tag_3),
    .io_out_tag_4(S8DP1_2_io_out_tag_4),
    .io_out_tag_5(S8DP1_2_io_out_tag_5),
    .io_out_tag_6(S8DP1_2_io_out_tag_6),
    .io_out_tag_7(S8DP1_2_io_out_tag_7),
    .io_result(S8DP1_2_io_result)
  );
  S8DP1 S8DP1_3( // @[STA_VDBB.scala 55:44:@8863.4]
    .clock(S8DP1_3_clock),
    .reset(S8DP1_3_reset),
    .io_int_in_A_0(S8DP1_3_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_3_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_3_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_3_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_3_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_3_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_3_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_3_io_int_in_A_7),
    .io_int_in_B(S8DP1_3_io_int_in_B),
    .io_tag_0(S8DP1_3_io_tag_0),
    .io_tag_1(S8DP1_3_io_tag_1),
    .io_tag_2(S8DP1_3_io_tag_2),
    .io_tag_3(S8DP1_3_io_tag_3),
    .io_tag_4(S8DP1_3_io_tag_4),
    .io_tag_5(S8DP1_3_io_tag_5),
    .io_tag_6(S8DP1_3_io_tag_6),
    .io_tag_7(S8DP1_3_io_tag_7),
    .io_out_tag_0(S8DP1_3_io_out_tag_0),
    .io_out_tag_1(S8DP1_3_io_out_tag_1),
    .io_out_tag_2(S8DP1_3_io_out_tag_2),
    .io_out_tag_3(S8DP1_3_io_out_tag_3),
    .io_out_tag_4(S8DP1_3_io_out_tag_4),
    .io_out_tag_5(S8DP1_3_io_out_tag_5),
    .io_out_tag_6(S8DP1_3_io_out_tag_6),
    .io_out_tag_7(S8DP1_3_io_out_tag_7),
    .io_result(S8DP1_3_io_result)
  );
  S8DP1 S8DP1_4( // @[STA_VDBB.scala 55:44:@8866.4]
    .clock(S8DP1_4_clock),
    .reset(S8DP1_4_reset),
    .io_int_in_A_0(S8DP1_4_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_4_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_4_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_4_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_4_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_4_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_4_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_4_io_int_in_A_7),
    .io_int_in_B(S8DP1_4_io_int_in_B),
    .io_tag_0(S8DP1_4_io_tag_0),
    .io_tag_1(S8DP1_4_io_tag_1),
    .io_tag_2(S8DP1_4_io_tag_2),
    .io_tag_3(S8DP1_4_io_tag_3),
    .io_tag_4(S8DP1_4_io_tag_4),
    .io_tag_5(S8DP1_4_io_tag_5),
    .io_tag_6(S8DP1_4_io_tag_6),
    .io_tag_7(S8DP1_4_io_tag_7),
    .io_out_tag_0(S8DP1_4_io_out_tag_0),
    .io_out_tag_1(S8DP1_4_io_out_tag_1),
    .io_out_tag_2(S8DP1_4_io_out_tag_2),
    .io_out_tag_3(S8DP1_4_io_out_tag_3),
    .io_out_tag_4(S8DP1_4_io_out_tag_4),
    .io_out_tag_5(S8DP1_4_io_out_tag_5),
    .io_out_tag_6(S8DP1_4_io_out_tag_6),
    .io_out_tag_7(S8DP1_4_io_out_tag_7),
    .io_result(S8DP1_4_io_result)
  );
  S8DP1 S8DP1_5( // @[STA_VDBB.scala 55:44:@8869.4]
    .clock(S8DP1_5_clock),
    .reset(S8DP1_5_reset),
    .io_int_in_A_0(S8DP1_5_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_5_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_5_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_5_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_5_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_5_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_5_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_5_io_int_in_A_7),
    .io_int_in_B(S8DP1_5_io_int_in_B),
    .io_tag_0(S8DP1_5_io_tag_0),
    .io_tag_1(S8DP1_5_io_tag_1),
    .io_tag_2(S8DP1_5_io_tag_2),
    .io_tag_3(S8DP1_5_io_tag_3),
    .io_tag_4(S8DP1_5_io_tag_4),
    .io_tag_5(S8DP1_5_io_tag_5),
    .io_tag_6(S8DP1_5_io_tag_6),
    .io_tag_7(S8DP1_5_io_tag_7),
    .io_out_tag_0(S8DP1_5_io_out_tag_0),
    .io_out_tag_1(S8DP1_5_io_out_tag_1),
    .io_out_tag_2(S8DP1_5_io_out_tag_2),
    .io_out_tag_3(S8DP1_5_io_out_tag_3),
    .io_out_tag_4(S8DP1_5_io_out_tag_4),
    .io_out_tag_5(S8DP1_5_io_out_tag_5),
    .io_out_tag_6(S8DP1_5_io_out_tag_6),
    .io_out_tag_7(S8DP1_5_io_out_tag_7),
    .io_result(S8DP1_5_io_result)
  );
  S8DP1 S8DP1_6( // @[STA_VDBB.scala 55:44:@8872.4]
    .clock(S8DP1_6_clock),
    .reset(S8DP1_6_reset),
    .io_int_in_A_0(S8DP1_6_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_6_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_6_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_6_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_6_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_6_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_6_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_6_io_int_in_A_7),
    .io_int_in_B(S8DP1_6_io_int_in_B),
    .io_tag_0(S8DP1_6_io_tag_0),
    .io_tag_1(S8DP1_6_io_tag_1),
    .io_tag_2(S8DP1_6_io_tag_2),
    .io_tag_3(S8DP1_6_io_tag_3),
    .io_tag_4(S8DP1_6_io_tag_4),
    .io_tag_5(S8DP1_6_io_tag_5),
    .io_tag_6(S8DP1_6_io_tag_6),
    .io_tag_7(S8DP1_6_io_tag_7),
    .io_out_tag_0(S8DP1_6_io_out_tag_0),
    .io_out_tag_1(S8DP1_6_io_out_tag_1),
    .io_out_tag_2(S8DP1_6_io_out_tag_2),
    .io_out_tag_3(S8DP1_6_io_out_tag_3),
    .io_out_tag_4(S8DP1_6_io_out_tag_4),
    .io_out_tag_5(S8DP1_6_io_out_tag_5),
    .io_out_tag_6(S8DP1_6_io_out_tag_6),
    .io_out_tag_7(S8DP1_6_io_out_tag_7),
    .io_result(S8DP1_6_io_result)
  );
  S8DP1 S8DP1_7( // @[STA_VDBB.scala 55:44:@8875.4]
    .clock(S8DP1_7_clock),
    .reset(S8DP1_7_reset),
    .io_int_in_A_0(S8DP1_7_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_7_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_7_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_7_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_7_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_7_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_7_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_7_io_int_in_A_7),
    .io_int_in_B(S8DP1_7_io_int_in_B),
    .io_tag_0(S8DP1_7_io_tag_0),
    .io_tag_1(S8DP1_7_io_tag_1),
    .io_tag_2(S8DP1_7_io_tag_2),
    .io_tag_3(S8DP1_7_io_tag_3),
    .io_tag_4(S8DP1_7_io_tag_4),
    .io_tag_5(S8DP1_7_io_tag_5),
    .io_tag_6(S8DP1_7_io_tag_6),
    .io_tag_7(S8DP1_7_io_tag_7),
    .io_out_tag_0(S8DP1_7_io_out_tag_0),
    .io_out_tag_1(S8DP1_7_io_out_tag_1),
    .io_out_tag_2(S8DP1_7_io_out_tag_2),
    .io_out_tag_3(S8DP1_7_io_out_tag_3),
    .io_out_tag_4(S8DP1_7_io_out_tag_4),
    .io_out_tag_5(S8DP1_7_io_out_tag_5),
    .io_out_tag_6(S8DP1_7_io_out_tag_6),
    .io_out_tag_7(S8DP1_7_io_out_tag_7),
    .io_result(S8DP1_7_io_result)
  );
  S8DP1 S8DP1_8( // @[STA_VDBB.scala 56:44:@9087.4]
    .clock(S8DP1_8_clock),
    .reset(S8DP1_8_reset),
    .io_int_in_A_0(S8DP1_8_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_8_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_8_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_8_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_8_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_8_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_8_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_8_io_int_in_A_7),
    .io_int_in_B(S8DP1_8_io_int_in_B),
    .io_tag_0(S8DP1_8_io_tag_0),
    .io_tag_1(S8DP1_8_io_tag_1),
    .io_tag_2(S8DP1_8_io_tag_2),
    .io_tag_3(S8DP1_8_io_tag_3),
    .io_tag_4(S8DP1_8_io_tag_4),
    .io_tag_5(S8DP1_8_io_tag_5),
    .io_tag_6(S8DP1_8_io_tag_6),
    .io_tag_7(S8DP1_8_io_tag_7),
    .io_out_tag_0(S8DP1_8_io_out_tag_0),
    .io_out_tag_1(S8DP1_8_io_out_tag_1),
    .io_out_tag_2(S8DP1_8_io_out_tag_2),
    .io_out_tag_3(S8DP1_8_io_out_tag_3),
    .io_out_tag_4(S8DP1_8_io_out_tag_4),
    .io_out_tag_5(S8DP1_8_io_out_tag_5),
    .io_out_tag_6(S8DP1_8_io_out_tag_6),
    .io_out_tag_7(S8DP1_8_io_out_tag_7),
    .io_result(S8DP1_8_io_result)
  );
  S8DP1 S8DP1_9( // @[STA_VDBB.scala 56:44:@9090.4]
    .clock(S8DP1_9_clock),
    .reset(S8DP1_9_reset),
    .io_int_in_A_0(S8DP1_9_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_9_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_9_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_9_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_9_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_9_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_9_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_9_io_int_in_A_7),
    .io_int_in_B(S8DP1_9_io_int_in_B),
    .io_tag_0(S8DP1_9_io_tag_0),
    .io_tag_1(S8DP1_9_io_tag_1),
    .io_tag_2(S8DP1_9_io_tag_2),
    .io_tag_3(S8DP1_9_io_tag_3),
    .io_tag_4(S8DP1_9_io_tag_4),
    .io_tag_5(S8DP1_9_io_tag_5),
    .io_tag_6(S8DP1_9_io_tag_6),
    .io_tag_7(S8DP1_9_io_tag_7),
    .io_out_tag_0(S8DP1_9_io_out_tag_0),
    .io_out_tag_1(S8DP1_9_io_out_tag_1),
    .io_out_tag_2(S8DP1_9_io_out_tag_2),
    .io_out_tag_3(S8DP1_9_io_out_tag_3),
    .io_out_tag_4(S8DP1_9_io_out_tag_4),
    .io_out_tag_5(S8DP1_9_io_out_tag_5),
    .io_out_tag_6(S8DP1_9_io_out_tag_6),
    .io_out_tag_7(S8DP1_9_io_out_tag_7),
    .io_result(S8DP1_9_io_result)
  );
  S8DP1 S8DP1_10( // @[STA_VDBB.scala 56:44:@9093.4]
    .clock(S8DP1_10_clock),
    .reset(S8DP1_10_reset),
    .io_int_in_A_0(S8DP1_10_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_10_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_10_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_10_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_10_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_10_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_10_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_10_io_int_in_A_7),
    .io_int_in_B(S8DP1_10_io_int_in_B),
    .io_tag_0(S8DP1_10_io_tag_0),
    .io_tag_1(S8DP1_10_io_tag_1),
    .io_tag_2(S8DP1_10_io_tag_2),
    .io_tag_3(S8DP1_10_io_tag_3),
    .io_tag_4(S8DP1_10_io_tag_4),
    .io_tag_5(S8DP1_10_io_tag_5),
    .io_tag_6(S8DP1_10_io_tag_6),
    .io_tag_7(S8DP1_10_io_tag_7),
    .io_out_tag_0(S8DP1_10_io_out_tag_0),
    .io_out_tag_1(S8DP1_10_io_out_tag_1),
    .io_out_tag_2(S8DP1_10_io_out_tag_2),
    .io_out_tag_3(S8DP1_10_io_out_tag_3),
    .io_out_tag_4(S8DP1_10_io_out_tag_4),
    .io_out_tag_5(S8DP1_10_io_out_tag_5),
    .io_out_tag_6(S8DP1_10_io_out_tag_6),
    .io_out_tag_7(S8DP1_10_io_out_tag_7),
    .io_result(S8DP1_10_io_result)
  );
  S8DP1 S8DP1_11( // @[STA_VDBB.scala 56:44:@9096.4]
    .clock(S8DP1_11_clock),
    .reset(S8DP1_11_reset),
    .io_int_in_A_0(S8DP1_11_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_11_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_11_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_11_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_11_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_11_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_11_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_11_io_int_in_A_7),
    .io_int_in_B(S8DP1_11_io_int_in_B),
    .io_tag_0(S8DP1_11_io_tag_0),
    .io_tag_1(S8DP1_11_io_tag_1),
    .io_tag_2(S8DP1_11_io_tag_2),
    .io_tag_3(S8DP1_11_io_tag_3),
    .io_tag_4(S8DP1_11_io_tag_4),
    .io_tag_5(S8DP1_11_io_tag_5),
    .io_tag_6(S8DP1_11_io_tag_6),
    .io_tag_7(S8DP1_11_io_tag_7),
    .io_out_tag_0(S8DP1_11_io_out_tag_0),
    .io_out_tag_1(S8DP1_11_io_out_tag_1),
    .io_out_tag_2(S8DP1_11_io_out_tag_2),
    .io_out_tag_3(S8DP1_11_io_out_tag_3),
    .io_out_tag_4(S8DP1_11_io_out_tag_4),
    .io_out_tag_5(S8DP1_11_io_out_tag_5),
    .io_out_tag_6(S8DP1_11_io_out_tag_6),
    .io_out_tag_7(S8DP1_11_io_out_tag_7),
    .io_result(S8DP1_11_io_result)
  );
  S8DP1 S8DP1_12( // @[STA_VDBB.scala 56:44:@9099.4]
    .clock(S8DP1_12_clock),
    .reset(S8DP1_12_reset),
    .io_int_in_A_0(S8DP1_12_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_12_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_12_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_12_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_12_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_12_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_12_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_12_io_int_in_A_7),
    .io_int_in_B(S8DP1_12_io_int_in_B),
    .io_tag_0(S8DP1_12_io_tag_0),
    .io_tag_1(S8DP1_12_io_tag_1),
    .io_tag_2(S8DP1_12_io_tag_2),
    .io_tag_3(S8DP1_12_io_tag_3),
    .io_tag_4(S8DP1_12_io_tag_4),
    .io_tag_5(S8DP1_12_io_tag_5),
    .io_tag_6(S8DP1_12_io_tag_6),
    .io_tag_7(S8DP1_12_io_tag_7),
    .io_out_tag_0(S8DP1_12_io_out_tag_0),
    .io_out_tag_1(S8DP1_12_io_out_tag_1),
    .io_out_tag_2(S8DP1_12_io_out_tag_2),
    .io_out_tag_3(S8DP1_12_io_out_tag_3),
    .io_out_tag_4(S8DP1_12_io_out_tag_4),
    .io_out_tag_5(S8DP1_12_io_out_tag_5),
    .io_out_tag_6(S8DP1_12_io_out_tag_6),
    .io_out_tag_7(S8DP1_12_io_out_tag_7),
    .io_result(S8DP1_12_io_result)
  );
  S8DP1 S8DP1_13( // @[STA_VDBB.scala 56:44:@9102.4]
    .clock(S8DP1_13_clock),
    .reset(S8DP1_13_reset),
    .io_int_in_A_0(S8DP1_13_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_13_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_13_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_13_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_13_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_13_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_13_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_13_io_int_in_A_7),
    .io_int_in_B(S8DP1_13_io_int_in_B),
    .io_tag_0(S8DP1_13_io_tag_0),
    .io_tag_1(S8DP1_13_io_tag_1),
    .io_tag_2(S8DP1_13_io_tag_2),
    .io_tag_3(S8DP1_13_io_tag_3),
    .io_tag_4(S8DP1_13_io_tag_4),
    .io_tag_5(S8DP1_13_io_tag_5),
    .io_tag_6(S8DP1_13_io_tag_6),
    .io_tag_7(S8DP1_13_io_tag_7),
    .io_out_tag_0(S8DP1_13_io_out_tag_0),
    .io_out_tag_1(S8DP1_13_io_out_tag_1),
    .io_out_tag_2(S8DP1_13_io_out_tag_2),
    .io_out_tag_3(S8DP1_13_io_out_tag_3),
    .io_out_tag_4(S8DP1_13_io_out_tag_4),
    .io_out_tag_5(S8DP1_13_io_out_tag_5),
    .io_out_tag_6(S8DP1_13_io_out_tag_6),
    .io_out_tag_7(S8DP1_13_io_out_tag_7),
    .io_result(S8DP1_13_io_result)
  );
  S8DP1 S8DP1_14( // @[STA_VDBB.scala 56:44:@9105.4]
    .clock(S8DP1_14_clock),
    .reset(S8DP1_14_reset),
    .io_int_in_A_0(S8DP1_14_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_14_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_14_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_14_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_14_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_14_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_14_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_14_io_int_in_A_7),
    .io_int_in_B(S8DP1_14_io_int_in_B),
    .io_tag_0(S8DP1_14_io_tag_0),
    .io_tag_1(S8DP1_14_io_tag_1),
    .io_tag_2(S8DP1_14_io_tag_2),
    .io_tag_3(S8DP1_14_io_tag_3),
    .io_tag_4(S8DP1_14_io_tag_4),
    .io_tag_5(S8DP1_14_io_tag_5),
    .io_tag_6(S8DP1_14_io_tag_6),
    .io_tag_7(S8DP1_14_io_tag_7),
    .io_out_tag_0(S8DP1_14_io_out_tag_0),
    .io_out_tag_1(S8DP1_14_io_out_tag_1),
    .io_out_tag_2(S8DP1_14_io_out_tag_2),
    .io_out_tag_3(S8DP1_14_io_out_tag_3),
    .io_out_tag_4(S8DP1_14_io_out_tag_4),
    .io_out_tag_5(S8DP1_14_io_out_tag_5),
    .io_out_tag_6(S8DP1_14_io_out_tag_6),
    .io_out_tag_7(S8DP1_14_io_out_tag_7),
    .io_result(S8DP1_14_io_result)
  );
  S8DP1 S8DP1_15( // @[STA_VDBB.scala 56:44:@9108.4]
    .clock(S8DP1_15_clock),
    .reset(S8DP1_15_reset),
    .io_int_in_A_0(S8DP1_15_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_15_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_15_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_15_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_15_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_15_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_15_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_15_io_int_in_A_7),
    .io_int_in_B(S8DP1_15_io_int_in_B),
    .io_tag_0(S8DP1_15_io_tag_0),
    .io_tag_1(S8DP1_15_io_tag_1),
    .io_tag_2(S8DP1_15_io_tag_2),
    .io_tag_3(S8DP1_15_io_tag_3),
    .io_tag_4(S8DP1_15_io_tag_4),
    .io_tag_5(S8DP1_15_io_tag_5),
    .io_tag_6(S8DP1_15_io_tag_6),
    .io_tag_7(S8DP1_15_io_tag_7),
    .io_out_tag_0(S8DP1_15_io_out_tag_0),
    .io_out_tag_1(S8DP1_15_io_out_tag_1),
    .io_out_tag_2(S8DP1_15_io_out_tag_2),
    .io_out_tag_3(S8DP1_15_io_out_tag_3),
    .io_out_tag_4(S8DP1_15_io_out_tag_4),
    .io_out_tag_5(S8DP1_15_io_out_tag_5),
    .io_out_tag_6(S8DP1_15_io_out_tag_6),
    .io_out_tag_7(S8DP1_15_io_out_tag_7),
    .io_result(S8DP1_15_io_result)
  );
  S8DP1 S8DP1_16( // @[STA_VDBB.scala 57:44:@9320.4]
    .clock(S8DP1_16_clock),
    .reset(S8DP1_16_reset),
    .io_int_in_A_0(S8DP1_16_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_16_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_16_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_16_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_16_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_16_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_16_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_16_io_int_in_A_7),
    .io_int_in_B(S8DP1_16_io_int_in_B),
    .io_tag_0(S8DP1_16_io_tag_0),
    .io_tag_1(S8DP1_16_io_tag_1),
    .io_tag_2(S8DP1_16_io_tag_2),
    .io_tag_3(S8DP1_16_io_tag_3),
    .io_tag_4(S8DP1_16_io_tag_4),
    .io_tag_5(S8DP1_16_io_tag_5),
    .io_tag_6(S8DP1_16_io_tag_6),
    .io_tag_7(S8DP1_16_io_tag_7),
    .io_out_tag_0(S8DP1_16_io_out_tag_0),
    .io_out_tag_1(S8DP1_16_io_out_tag_1),
    .io_out_tag_2(S8DP1_16_io_out_tag_2),
    .io_out_tag_3(S8DP1_16_io_out_tag_3),
    .io_out_tag_4(S8DP1_16_io_out_tag_4),
    .io_out_tag_5(S8DP1_16_io_out_tag_5),
    .io_out_tag_6(S8DP1_16_io_out_tag_6),
    .io_out_tag_7(S8DP1_16_io_out_tag_7),
    .io_result(S8DP1_16_io_result)
  );
  S8DP1 S8DP1_17( // @[STA_VDBB.scala 57:44:@9323.4]
    .clock(S8DP1_17_clock),
    .reset(S8DP1_17_reset),
    .io_int_in_A_0(S8DP1_17_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_17_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_17_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_17_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_17_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_17_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_17_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_17_io_int_in_A_7),
    .io_int_in_B(S8DP1_17_io_int_in_B),
    .io_tag_0(S8DP1_17_io_tag_0),
    .io_tag_1(S8DP1_17_io_tag_1),
    .io_tag_2(S8DP1_17_io_tag_2),
    .io_tag_3(S8DP1_17_io_tag_3),
    .io_tag_4(S8DP1_17_io_tag_4),
    .io_tag_5(S8DP1_17_io_tag_5),
    .io_tag_6(S8DP1_17_io_tag_6),
    .io_tag_7(S8DP1_17_io_tag_7),
    .io_out_tag_0(S8DP1_17_io_out_tag_0),
    .io_out_tag_1(S8DP1_17_io_out_tag_1),
    .io_out_tag_2(S8DP1_17_io_out_tag_2),
    .io_out_tag_3(S8DP1_17_io_out_tag_3),
    .io_out_tag_4(S8DP1_17_io_out_tag_4),
    .io_out_tag_5(S8DP1_17_io_out_tag_5),
    .io_out_tag_6(S8DP1_17_io_out_tag_6),
    .io_out_tag_7(S8DP1_17_io_out_tag_7),
    .io_result(S8DP1_17_io_result)
  );
  S8DP1 S8DP1_18( // @[STA_VDBB.scala 57:44:@9326.4]
    .clock(S8DP1_18_clock),
    .reset(S8DP1_18_reset),
    .io_int_in_A_0(S8DP1_18_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_18_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_18_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_18_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_18_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_18_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_18_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_18_io_int_in_A_7),
    .io_int_in_B(S8DP1_18_io_int_in_B),
    .io_tag_0(S8DP1_18_io_tag_0),
    .io_tag_1(S8DP1_18_io_tag_1),
    .io_tag_2(S8DP1_18_io_tag_2),
    .io_tag_3(S8DP1_18_io_tag_3),
    .io_tag_4(S8DP1_18_io_tag_4),
    .io_tag_5(S8DP1_18_io_tag_5),
    .io_tag_6(S8DP1_18_io_tag_6),
    .io_tag_7(S8DP1_18_io_tag_7),
    .io_out_tag_0(S8DP1_18_io_out_tag_0),
    .io_out_tag_1(S8DP1_18_io_out_tag_1),
    .io_out_tag_2(S8DP1_18_io_out_tag_2),
    .io_out_tag_3(S8DP1_18_io_out_tag_3),
    .io_out_tag_4(S8DP1_18_io_out_tag_4),
    .io_out_tag_5(S8DP1_18_io_out_tag_5),
    .io_out_tag_6(S8DP1_18_io_out_tag_6),
    .io_out_tag_7(S8DP1_18_io_out_tag_7),
    .io_result(S8DP1_18_io_result)
  );
  S8DP1 S8DP1_19( // @[STA_VDBB.scala 57:44:@9329.4]
    .clock(S8DP1_19_clock),
    .reset(S8DP1_19_reset),
    .io_int_in_A_0(S8DP1_19_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_19_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_19_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_19_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_19_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_19_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_19_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_19_io_int_in_A_7),
    .io_int_in_B(S8DP1_19_io_int_in_B),
    .io_tag_0(S8DP1_19_io_tag_0),
    .io_tag_1(S8DP1_19_io_tag_1),
    .io_tag_2(S8DP1_19_io_tag_2),
    .io_tag_3(S8DP1_19_io_tag_3),
    .io_tag_4(S8DP1_19_io_tag_4),
    .io_tag_5(S8DP1_19_io_tag_5),
    .io_tag_6(S8DP1_19_io_tag_6),
    .io_tag_7(S8DP1_19_io_tag_7),
    .io_out_tag_0(S8DP1_19_io_out_tag_0),
    .io_out_tag_1(S8DP1_19_io_out_tag_1),
    .io_out_tag_2(S8DP1_19_io_out_tag_2),
    .io_out_tag_3(S8DP1_19_io_out_tag_3),
    .io_out_tag_4(S8DP1_19_io_out_tag_4),
    .io_out_tag_5(S8DP1_19_io_out_tag_5),
    .io_out_tag_6(S8DP1_19_io_out_tag_6),
    .io_out_tag_7(S8DP1_19_io_out_tag_7),
    .io_result(S8DP1_19_io_result)
  );
  S8DP1 S8DP1_20( // @[STA_VDBB.scala 57:44:@9332.4]
    .clock(S8DP1_20_clock),
    .reset(S8DP1_20_reset),
    .io_int_in_A_0(S8DP1_20_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_20_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_20_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_20_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_20_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_20_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_20_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_20_io_int_in_A_7),
    .io_int_in_B(S8DP1_20_io_int_in_B),
    .io_tag_0(S8DP1_20_io_tag_0),
    .io_tag_1(S8DP1_20_io_tag_1),
    .io_tag_2(S8DP1_20_io_tag_2),
    .io_tag_3(S8DP1_20_io_tag_3),
    .io_tag_4(S8DP1_20_io_tag_4),
    .io_tag_5(S8DP1_20_io_tag_5),
    .io_tag_6(S8DP1_20_io_tag_6),
    .io_tag_7(S8DP1_20_io_tag_7),
    .io_out_tag_0(S8DP1_20_io_out_tag_0),
    .io_out_tag_1(S8DP1_20_io_out_tag_1),
    .io_out_tag_2(S8DP1_20_io_out_tag_2),
    .io_out_tag_3(S8DP1_20_io_out_tag_3),
    .io_out_tag_4(S8DP1_20_io_out_tag_4),
    .io_out_tag_5(S8DP1_20_io_out_tag_5),
    .io_out_tag_6(S8DP1_20_io_out_tag_6),
    .io_out_tag_7(S8DP1_20_io_out_tag_7),
    .io_result(S8DP1_20_io_result)
  );
  S8DP1 S8DP1_21( // @[STA_VDBB.scala 57:44:@9335.4]
    .clock(S8DP1_21_clock),
    .reset(S8DP1_21_reset),
    .io_int_in_A_0(S8DP1_21_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_21_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_21_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_21_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_21_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_21_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_21_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_21_io_int_in_A_7),
    .io_int_in_B(S8DP1_21_io_int_in_B),
    .io_tag_0(S8DP1_21_io_tag_0),
    .io_tag_1(S8DP1_21_io_tag_1),
    .io_tag_2(S8DP1_21_io_tag_2),
    .io_tag_3(S8DP1_21_io_tag_3),
    .io_tag_4(S8DP1_21_io_tag_4),
    .io_tag_5(S8DP1_21_io_tag_5),
    .io_tag_6(S8DP1_21_io_tag_6),
    .io_tag_7(S8DP1_21_io_tag_7),
    .io_out_tag_0(S8DP1_21_io_out_tag_0),
    .io_out_tag_1(S8DP1_21_io_out_tag_1),
    .io_out_tag_2(S8DP1_21_io_out_tag_2),
    .io_out_tag_3(S8DP1_21_io_out_tag_3),
    .io_out_tag_4(S8DP1_21_io_out_tag_4),
    .io_out_tag_5(S8DP1_21_io_out_tag_5),
    .io_out_tag_6(S8DP1_21_io_out_tag_6),
    .io_out_tag_7(S8DP1_21_io_out_tag_7),
    .io_result(S8DP1_21_io_result)
  );
  S8DP1 S8DP1_22( // @[STA_VDBB.scala 57:44:@9338.4]
    .clock(S8DP1_22_clock),
    .reset(S8DP1_22_reset),
    .io_int_in_A_0(S8DP1_22_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_22_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_22_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_22_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_22_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_22_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_22_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_22_io_int_in_A_7),
    .io_int_in_B(S8DP1_22_io_int_in_B),
    .io_tag_0(S8DP1_22_io_tag_0),
    .io_tag_1(S8DP1_22_io_tag_1),
    .io_tag_2(S8DP1_22_io_tag_2),
    .io_tag_3(S8DP1_22_io_tag_3),
    .io_tag_4(S8DP1_22_io_tag_4),
    .io_tag_5(S8DP1_22_io_tag_5),
    .io_tag_6(S8DP1_22_io_tag_6),
    .io_tag_7(S8DP1_22_io_tag_7),
    .io_out_tag_0(S8DP1_22_io_out_tag_0),
    .io_out_tag_1(S8DP1_22_io_out_tag_1),
    .io_out_tag_2(S8DP1_22_io_out_tag_2),
    .io_out_tag_3(S8DP1_22_io_out_tag_3),
    .io_out_tag_4(S8DP1_22_io_out_tag_4),
    .io_out_tag_5(S8DP1_22_io_out_tag_5),
    .io_out_tag_6(S8DP1_22_io_out_tag_6),
    .io_out_tag_7(S8DP1_22_io_out_tag_7),
    .io_result(S8DP1_22_io_result)
  );
  S8DP1 S8DP1_23( // @[STA_VDBB.scala 57:44:@9341.4]
    .clock(S8DP1_23_clock),
    .reset(S8DP1_23_reset),
    .io_int_in_A_0(S8DP1_23_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_23_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_23_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_23_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_23_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_23_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_23_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_23_io_int_in_A_7),
    .io_int_in_B(S8DP1_23_io_int_in_B),
    .io_tag_0(S8DP1_23_io_tag_0),
    .io_tag_1(S8DP1_23_io_tag_1),
    .io_tag_2(S8DP1_23_io_tag_2),
    .io_tag_3(S8DP1_23_io_tag_3),
    .io_tag_4(S8DP1_23_io_tag_4),
    .io_tag_5(S8DP1_23_io_tag_5),
    .io_tag_6(S8DP1_23_io_tag_6),
    .io_tag_7(S8DP1_23_io_tag_7),
    .io_out_tag_0(S8DP1_23_io_out_tag_0),
    .io_out_tag_1(S8DP1_23_io_out_tag_1),
    .io_out_tag_2(S8DP1_23_io_out_tag_2),
    .io_out_tag_3(S8DP1_23_io_out_tag_3),
    .io_out_tag_4(S8DP1_23_io_out_tag_4),
    .io_out_tag_5(S8DP1_23_io_out_tag_5),
    .io_out_tag_6(S8DP1_23_io_out_tag_6),
    .io_out_tag_7(S8DP1_23_io_out_tag_7),
    .io_result(S8DP1_23_io_result)
  );
  S8DP1 S8DP1_24( // @[STA_VDBB.scala 58:44:@9553.4]
    .clock(S8DP1_24_clock),
    .reset(S8DP1_24_reset),
    .io_int_in_A_0(S8DP1_24_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_24_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_24_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_24_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_24_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_24_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_24_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_24_io_int_in_A_7),
    .io_int_in_B(S8DP1_24_io_int_in_B),
    .io_tag_0(S8DP1_24_io_tag_0),
    .io_tag_1(S8DP1_24_io_tag_1),
    .io_tag_2(S8DP1_24_io_tag_2),
    .io_tag_3(S8DP1_24_io_tag_3),
    .io_tag_4(S8DP1_24_io_tag_4),
    .io_tag_5(S8DP1_24_io_tag_5),
    .io_tag_6(S8DP1_24_io_tag_6),
    .io_tag_7(S8DP1_24_io_tag_7),
    .io_out_tag_0(S8DP1_24_io_out_tag_0),
    .io_out_tag_1(S8DP1_24_io_out_tag_1),
    .io_out_tag_2(S8DP1_24_io_out_tag_2),
    .io_out_tag_3(S8DP1_24_io_out_tag_3),
    .io_out_tag_4(S8DP1_24_io_out_tag_4),
    .io_out_tag_5(S8DP1_24_io_out_tag_5),
    .io_out_tag_6(S8DP1_24_io_out_tag_6),
    .io_out_tag_7(S8DP1_24_io_out_tag_7),
    .io_result(S8DP1_24_io_result)
  );
  S8DP1 S8DP1_25( // @[STA_VDBB.scala 58:44:@9556.4]
    .clock(S8DP1_25_clock),
    .reset(S8DP1_25_reset),
    .io_int_in_A_0(S8DP1_25_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_25_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_25_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_25_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_25_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_25_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_25_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_25_io_int_in_A_7),
    .io_int_in_B(S8DP1_25_io_int_in_B),
    .io_tag_0(S8DP1_25_io_tag_0),
    .io_tag_1(S8DP1_25_io_tag_1),
    .io_tag_2(S8DP1_25_io_tag_2),
    .io_tag_3(S8DP1_25_io_tag_3),
    .io_tag_4(S8DP1_25_io_tag_4),
    .io_tag_5(S8DP1_25_io_tag_5),
    .io_tag_6(S8DP1_25_io_tag_6),
    .io_tag_7(S8DP1_25_io_tag_7),
    .io_out_tag_0(S8DP1_25_io_out_tag_0),
    .io_out_tag_1(S8DP1_25_io_out_tag_1),
    .io_out_tag_2(S8DP1_25_io_out_tag_2),
    .io_out_tag_3(S8DP1_25_io_out_tag_3),
    .io_out_tag_4(S8DP1_25_io_out_tag_4),
    .io_out_tag_5(S8DP1_25_io_out_tag_5),
    .io_out_tag_6(S8DP1_25_io_out_tag_6),
    .io_out_tag_7(S8DP1_25_io_out_tag_7),
    .io_result(S8DP1_25_io_result)
  );
  S8DP1 S8DP1_26( // @[STA_VDBB.scala 58:44:@9559.4]
    .clock(S8DP1_26_clock),
    .reset(S8DP1_26_reset),
    .io_int_in_A_0(S8DP1_26_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_26_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_26_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_26_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_26_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_26_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_26_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_26_io_int_in_A_7),
    .io_int_in_B(S8DP1_26_io_int_in_B),
    .io_tag_0(S8DP1_26_io_tag_0),
    .io_tag_1(S8DP1_26_io_tag_1),
    .io_tag_2(S8DP1_26_io_tag_2),
    .io_tag_3(S8DP1_26_io_tag_3),
    .io_tag_4(S8DP1_26_io_tag_4),
    .io_tag_5(S8DP1_26_io_tag_5),
    .io_tag_6(S8DP1_26_io_tag_6),
    .io_tag_7(S8DP1_26_io_tag_7),
    .io_out_tag_0(S8DP1_26_io_out_tag_0),
    .io_out_tag_1(S8DP1_26_io_out_tag_1),
    .io_out_tag_2(S8DP1_26_io_out_tag_2),
    .io_out_tag_3(S8DP1_26_io_out_tag_3),
    .io_out_tag_4(S8DP1_26_io_out_tag_4),
    .io_out_tag_5(S8DP1_26_io_out_tag_5),
    .io_out_tag_6(S8DP1_26_io_out_tag_6),
    .io_out_tag_7(S8DP1_26_io_out_tag_7),
    .io_result(S8DP1_26_io_result)
  );
  S8DP1 S8DP1_27( // @[STA_VDBB.scala 58:44:@9562.4]
    .clock(S8DP1_27_clock),
    .reset(S8DP1_27_reset),
    .io_int_in_A_0(S8DP1_27_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_27_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_27_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_27_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_27_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_27_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_27_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_27_io_int_in_A_7),
    .io_int_in_B(S8DP1_27_io_int_in_B),
    .io_tag_0(S8DP1_27_io_tag_0),
    .io_tag_1(S8DP1_27_io_tag_1),
    .io_tag_2(S8DP1_27_io_tag_2),
    .io_tag_3(S8DP1_27_io_tag_3),
    .io_tag_4(S8DP1_27_io_tag_4),
    .io_tag_5(S8DP1_27_io_tag_5),
    .io_tag_6(S8DP1_27_io_tag_6),
    .io_tag_7(S8DP1_27_io_tag_7),
    .io_out_tag_0(S8DP1_27_io_out_tag_0),
    .io_out_tag_1(S8DP1_27_io_out_tag_1),
    .io_out_tag_2(S8DP1_27_io_out_tag_2),
    .io_out_tag_3(S8DP1_27_io_out_tag_3),
    .io_out_tag_4(S8DP1_27_io_out_tag_4),
    .io_out_tag_5(S8DP1_27_io_out_tag_5),
    .io_out_tag_6(S8DP1_27_io_out_tag_6),
    .io_out_tag_7(S8DP1_27_io_out_tag_7),
    .io_result(S8DP1_27_io_result)
  );
  S8DP1 S8DP1_28( // @[STA_VDBB.scala 58:44:@9565.4]
    .clock(S8DP1_28_clock),
    .reset(S8DP1_28_reset),
    .io_int_in_A_0(S8DP1_28_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_28_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_28_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_28_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_28_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_28_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_28_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_28_io_int_in_A_7),
    .io_int_in_B(S8DP1_28_io_int_in_B),
    .io_tag_0(S8DP1_28_io_tag_0),
    .io_tag_1(S8DP1_28_io_tag_1),
    .io_tag_2(S8DP1_28_io_tag_2),
    .io_tag_3(S8DP1_28_io_tag_3),
    .io_tag_4(S8DP1_28_io_tag_4),
    .io_tag_5(S8DP1_28_io_tag_5),
    .io_tag_6(S8DP1_28_io_tag_6),
    .io_tag_7(S8DP1_28_io_tag_7),
    .io_out_tag_0(S8DP1_28_io_out_tag_0),
    .io_out_tag_1(S8DP1_28_io_out_tag_1),
    .io_out_tag_2(S8DP1_28_io_out_tag_2),
    .io_out_tag_3(S8DP1_28_io_out_tag_3),
    .io_out_tag_4(S8DP1_28_io_out_tag_4),
    .io_out_tag_5(S8DP1_28_io_out_tag_5),
    .io_out_tag_6(S8DP1_28_io_out_tag_6),
    .io_out_tag_7(S8DP1_28_io_out_tag_7),
    .io_result(S8DP1_28_io_result)
  );
  S8DP1 S8DP1_29( // @[STA_VDBB.scala 58:44:@9568.4]
    .clock(S8DP1_29_clock),
    .reset(S8DP1_29_reset),
    .io_int_in_A_0(S8DP1_29_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_29_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_29_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_29_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_29_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_29_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_29_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_29_io_int_in_A_7),
    .io_int_in_B(S8DP1_29_io_int_in_B),
    .io_tag_0(S8DP1_29_io_tag_0),
    .io_tag_1(S8DP1_29_io_tag_1),
    .io_tag_2(S8DP1_29_io_tag_2),
    .io_tag_3(S8DP1_29_io_tag_3),
    .io_tag_4(S8DP1_29_io_tag_4),
    .io_tag_5(S8DP1_29_io_tag_5),
    .io_tag_6(S8DP1_29_io_tag_6),
    .io_tag_7(S8DP1_29_io_tag_7),
    .io_out_tag_0(S8DP1_29_io_out_tag_0),
    .io_out_tag_1(S8DP1_29_io_out_tag_1),
    .io_out_tag_2(S8DP1_29_io_out_tag_2),
    .io_out_tag_3(S8DP1_29_io_out_tag_3),
    .io_out_tag_4(S8DP1_29_io_out_tag_4),
    .io_out_tag_5(S8DP1_29_io_out_tag_5),
    .io_out_tag_6(S8DP1_29_io_out_tag_6),
    .io_out_tag_7(S8DP1_29_io_out_tag_7),
    .io_result(S8DP1_29_io_result)
  );
  S8DP1 S8DP1_30( // @[STA_VDBB.scala 58:44:@9571.4]
    .clock(S8DP1_30_clock),
    .reset(S8DP1_30_reset),
    .io_int_in_A_0(S8DP1_30_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_30_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_30_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_30_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_30_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_30_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_30_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_30_io_int_in_A_7),
    .io_int_in_B(S8DP1_30_io_int_in_B),
    .io_tag_0(S8DP1_30_io_tag_0),
    .io_tag_1(S8DP1_30_io_tag_1),
    .io_tag_2(S8DP1_30_io_tag_2),
    .io_tag_3(S8DP1_30_io_tag_3),
    .io_tag_4(S8DP1_30_io_tag_4),
    .io_tag_5(S8DP1_30_io_tag_5),
    .io_tag_6(S8DP1_30_io_tag_6),
    .io_tag_7(S8DP1_30_io_tag_7),
    .io_out_tag_0(S8DP1_30_io_out_tag_0),
    .io_out_tag_1(S8DP1_30_io_out_tag_1),
    .io_out_tag_2(S8DP1_30_io_out_tag_2),
    .io_out_tag_3(S8DP1_30_io_out_tag_3),
    .io_out_tag_4(S8DP1_30_io_out_tag_4),
    .io_out_tag_5(S8DP1_30_io_out_tag_5),
    .io_out_tag_6(S8DP1_30_io_out_tag_6),
    .io_out_tag_7(S8DP1_30_io_out_tag_7),
    .io_result(S8DP1_30_io_result)
  );
  S8DP1 S8DP1_31( // @[STA_VDBB.scala 58:44:@9574.4]
    .clock(S8DP1_31_clock),
    .reset(S8DP1_31_reset),
    .io_int_in_A_0(S8DP1_31_io_int_in_A_0),
    .io_int_in_A_1(S8DP1_31_io_int_in_A_1),
    .io_int_in_A_2(S8DP1_31_io_int_in_A_2),
    .io_int_in_A_3(S8DP1_31_io_int_in_A_3),
    .io_int_in_A_4(S8DP1_31_io_int_in_A_4),
    .io_int_in_A_5(S8DP1_31_io_int_in_A_5),
    .io_int_in_A_6(S8DP1_31_io_int_in_A_6),
    .io_int_in_A_7(S8DP1_31_io_int_in_A_7),
    .io_int_in_B(S8DP1_31_io_int_in_B),
    .io_tag_0(S8DP1_31_io_tag_0),
    .io_tag_1(S8DP1_31_io_tag_1),
    .io_tag_2(S8DP1_31_io_tag_2),
    .io_tag_3(S8DP1_31_io_tag_3),
    .io_tag_4(S8DP1_31_io_tag_4),
    .io_tag_5(S8DP1_31_io_tag_5),
    .io_tag_6(S8DP1_31_io_tag_6),
    .io_tag_7(S8DP1_31_io_tag_7),
    .io_out_tag_0(S8DP1_31_io_out_tag_0),
    .io_out_tag_1(S8DP1_31_io_out_tag_1),
    .io_out_tag_2(S8DP1_31_io_out_tag_2),
    .io_out_tag_3(S8DP1_31_io_out_tag_3),
    .io_out_tag_4(S8DP1_31_io_out_tag_4),
    .io_out_tag_5(S8DP1_31_io_out_tag_5),
    .io_out_tag_6(S8DP1_31_io_out_tag_6),
    .io_out_tag_7(S8DP1_31_io_out_tag_7),
    .io_result(S8DP1_31_io_result)
  );
  FF4 ffb1( // @[STA_VDBB.scala 68:20:@9786.4]
    .clock(ffb1_clock),
    .reset(ffb1_reset),
    .io_in_data_0_0(ffb1_io_in_data_0_0),
    .io_in_data_0_1(ffb1_io_in_data_0_1),
    .io_in_data_0_2(ffb1_io_in_data_0_2),
    .io_in_data_0_3(ffb1_io_in_data_0_3),
    .io_in_data_0_4(ffb1_io_in_data_0_4),
    .io_in_data_0_5(ffb1_io_in_data_0_5),
    .io_in_data_0_6(ffb1_io_in_data_0_6),
    .io_in_data_0_7(ffb1_io_in_data_0_7),
    .io_in_data_1_0(ffb1_io_in_data_1_0),
    .io_in_data_1_1(ffb1_io_in_data_1_1),
    .io_in_data_1_2(ffb1_io_in_data_1_2),
    .io_in_data_1_3(ffb1_io_in_data_1_3),
    .io_in_data_1_4(ffb1_io_in_data_1_4),
    .io_in_data_1_5(ffb1_io_in_data_1_5),
    .io_in_data_1_6(ffb1_io_in_data_1_6),
    .io_in_data_1_7(ffb1_io_in_data_1_7),
    .io_in_data_2_0(ffb1_io_in_data_2_0),
    .io_in_data_2_1(ffb1_io_in_data_2_1),
    .io_in_data_2_2(ffb1_io_in_data_2_2),
    .io_in_data_2_3(ffb1_io_in_data_2_3),
    .io_in_data_2_4(ffb1_io_in_data_2_4),
    .io_in_data_2_5(ffb1_io_in_data_2_5),
    .io_in_data_2_6(ffb1_io_in_data_2_6),
    .io_in_data_2_7(ffb1_io_in_data_2_7),
    .io_in_data_3_0(ffb1_io_in_data_3_0),
    .io_in_data_3_1(ffb1_io_in_data_3_1),
    .io_in_data_3_2(ffb1_io_in_data_3_2),
    .io_in_data_3_3(ffb1_io_in_data_3_3),
    .io_in_data_3_4(ffb1_io_in_data_3_4),
    .io_in_data_3_5(ffb1_io_in_data_3_5),
    .io_in_data_3_6(ffb1_io_in_data_3_6),
    .io_in_data_3_7(ffb1_io_in_data_3_7),
    .io_in_tag_0_0(ffb1_io_in_tag_0_0),
    .io_in_tag_0_1(ffb1_io_in_tag_0_1),
    .io_in_tag_0_2(ffb1_io_in_tag_0_2),
    .io_in_tag_0_3(ffb1_io_in_tag_0_3),
    .io_in_tag_0_4(ffb1_io_in_tag_0_4),
    .io_in_tag_0_5(ffb1_io_in_tag_0_5),
    .io_in_tag_0_6(ffb1_io_in_tag_0_6),
    .io_in_tag_0_7(ffb1_io_in_tag_0_7),
    .io_in_tag_1_0(ffb1_io_in_tag_1_0),
    .io_in_tag_1_1(ffb1_io_in_tag_1_1),
    .io_in_tag_1_2(ffb1_io_in_tag_1_2),
    .io_in_tag_1_3(ffb1_io_in_tag_1_3),
    .io_in_tag_1_4(ffb1_io_in_tag_1_4),
    .io_in_tag_1_5(ffb1_io_in_tag_1_5),
    .io_in_tag_1_6(ffb1_io_in_tag_1_6),
    .io_in_tag_1_7(ffb1_io_in_tag_1_7),
    .io_in_tag_2_0(ffb1_io_in_tag_2_0),
    .io_in_tag_2_1(ffb1_io_in_tag_2_1),
    .io_in_tag_2_2(ffb1_io_in_tag_2_2),
    .io_in_tag_2_3(ffb1_io_in_tag_2_3),
    .io_in_tag_2_4(ffb1_io_in_tag_2_4),
    .io_in_tag_2_5(ffb1_io_in_tag_2_5),
    .io_in_tag_2_6(ffb1_io_in_tag_2_6),
    .io_in_tag_2_7(ffb1_io_in_tag_2_7),
    .io_in_tag_3_0(ffb1_io_in_tag_3_0),
    .io_in_tag_3_1(ffb1_io_in_tag_3_1),
    .io_in_tag_3_2(ffb1_io_in_tag_3_2),
    .io_in_tag_3_3(ffb1_io_in_tag_3_3),
    .io_in_tag_3_4(ffb1_io_in_tag_3_4),
    .io_in_tag_3_5(ffb1_io_in_tag_3_5),
    .io_in_tag_3_6(ffb1_io_in_tag_3_6),
    .io_in_tag_3_7(ffb1_io_in_tag_3_7),
    .io_out_data_0_0(ffb1_io_out_data_0_0),
    .io_out_data_0_1(ffb1_io_out_data_0_1),
    .io_out_data_0_2(ffb1_io_out_data_0_2),
    .io_out_data_0_3(ffb1_io_out_data_0_3),
    .io_out_data_0_4(ffb1_io_out_data_0_4),
    .io_out_data_0_5(ffb1_io_out_data_0_5),
    .io_out_data_0_6(ffb1_io_out_data_0_6),
    .io_out_data_0_7(ffb1_io_out_data_0_7),
    .io_out_data_1_0(ffb1_io_out_data_1_0),
    .io_out_data_1_1(ffb1_io_out_data_1_1),
    .io_out_data_1_2(ffb1_io_out_data_1_2),
    .io_out_data_1_3(ffb1_io_out_data_1_3),
    .io_out_data_1_4(ffb1_io_out_data_1_4),
    .io_out_data_1_5(ffb1_io_out_data_1_5),
    .io_out_data_1_6(ffb1_io_out_data_1_6),
    .io_out_data_1_7(ffb1_io_out_data_1_7),
    .io_out_data_2_0(ffb1_io_out_data_2_0),
    .io_out_data_2_1(ffb1_io_out_data_2_1),
    .io_out_data_2_2(ffb1_io_out_data_2_2),
    .io_out_data_2_3(ffb1_io_out_data_2_3),
    .io_out_data_2_4(ffb1_io_out_data_2_4),
    .io_out_data_2_5(ffb1_io_out_data_2_5),
    .io_out_data_2_6(ffb1_io_out_data_2_6),
    .io_out_data_2_7(ffb1_io_out_data_2_7),
    .io_out_data_3_0(ffb1_io_out_data_3_0),
    .io_out_data_3_1(ffb1_io_out_data_3_1),
    .io_out_data_3_2(ffb1_io_out_data_3_2),
    .io_out_data_3_3(ffb1_io_out_data_3_3),
    .io_out_data_3_4(ffb1_io_out_data_3_4),
    .io_out_data_3_5(ffb1_io_out_data_3_5),
    .io_out_data_3_6(ffb1_io_out_data_3_6),
    .io_out_data_3_7(ffb1_io_out_data_3_7),
    .io_out_tag_0_0(ffb1_io_out_tag_0_0),
    .io_out_tag_0_1(ffb1_io_out_tag_0_1),
    .io_out_tag_0_2(ffb1_io_out_tag_0_2),
    .io_out_tag_0_3(ffb1_io_out_tag_0_3),
    .io_out_tag_0_4(ffb1_io_out_tag_0_4),
    .io_out_tag_0_5(ffb1_io_out_tag_0_5),
    .io_out_tag_0_6(ffb1_io_out_tag_0_6),
    .io_out_tag_0_7(ffb1_io_out_tag_0_7),
    .io_out_tag_1_0(ffb1_io_out_tag_1_0),
    .io_out_tag_1_1(ffb1_io_out_tag_1_1),
    .io_out_tag_1_2(ffb1_io_out_tag_1_2),
    .io_out_tag_1_3(ffb1_io_out_tag_1_3),
    .io_out_tag_1_4(ffb1_io_out_tag_1_4),
    .io_out_tag_1_5(ffb1_io_out_tag_1_5),
    .io_out_tag_1_6(ffb1_io_out_tag_1_6),
    .io_out_tag_1_7(ffb1_io_out_tag_1_7),
    .io_out_tag_2_0(ffb1_io_out_tag_2_0),
    .io_out_tag_2_1(ffb1_io_out_tag_2_1),
    .io_out_tag_2_2(ffb1_io_out_tag_2_2),
    .io_out_tag_2_3(ffb1_io_out_tag_2_3),
    .io_out_tag_2_4(ffb1_io_out_tag_2_4),
    .io_out_tag_2_5(ffb1_io_out_tag_2_5),
    .io_out_tag_2_6(ffb1_io_out_tag_2_6),
    .io_out_tag_2_7(ffb1_io_out_tag_2_7),
    .io_out_tag_3_0(ffb1_io_out_tag_3_0),
    .io_out_tag_3_1(ffb1_io_out_tag_3_1),
    .io_out_tag_3_2(ffb1_io_out_tag_3_2),
    .io_out_tag_3_3(ffb1_io_out_tag_3_3),
    .io_out_tag_3_4(ffb1_io_out_tag_3_4),
    .io_out_tag_3_5(ffb1_io_out_tag_3_5),
    .io_out_tag_3_6(ffb1_io_out_tag_3_6),
    .io_out_tag_3_7(ffb1_io_out_tag_3_7)
  );
  FF4 ffb2( // @[STA_VDBB.scala 69:20:@9789.4]
    .clock(ffb2_clock),
    .reset(ffb2_reset),
    .io_in_data_0_0(ffb2_io_in_data_0_0),
    .io_in_data_0_1(ffb2_io_in_data_0_1),
    .io_in_data_0_2(ffb2_io_in_data_0_2),
    .io_in_data_0_3(ffb2_io_in_data_0_3),
    .io_in_data_0_4(ffb2_io_in_data_0_4),
    .io_in_data_0_5(ffb2_io_in_data_0_5),
    .io_in_data_0_6(ffb2_io_in_data_0_6),
    .io_in_data_0_7(ffb2_io_in_data_0_7),
    .io_in_data_1_0(ffb2_io_in_data_1_0),
    .io_in_data_1_1(ffb2_io_in_data_1_1),
    .io_in_data_1_2(ffb2_io_in_data_1_2),
    .io_in_data_1_3(ffb2_io_in_data_1_3),
    .io_in_data_1_4(ffb2_io_in_data_1_4),
    .io_in_data_1_5(ffb2_io_in_data_1_5),
    .io_in_data_1_6(ffb2_io_in_data_1_6),
    .io_in_data_1_7(ffb2_io_in_data_1_7),
    .io_in_data_2_0(ffb2_io_in_data_2_0),
    .io_in_data_2_1(ffb2_io_in_data_2_1),
    .io_in_data_2_2(ffb2_io_in_data_2_2),
    .io_in_data_2_3(ffb2_io_in_data_2_3),
    .io_in_data_2_4(ffb2_io_in_data_2_4),
    .io_in_data_2_5(ffb2_io_in_data_2_5),
    .io_in_data_2_6(ffb2_io_in_data_2_6),
    .io_in_data_2_7(ffb2_io_in_data_2_7),
    .io_in_data_3_0(ffb2_io_in_data_3_0),
    .io_in_data_3_1(ffb2_io_in_data_3_1),
    .io_in_data_3_2(ffb2_io_in_data_3_2),
    .io_in_data_3_3(ffb2_io_in_data_3_3),
    .io_in_data_3_4(ffb2_io_in_data_3_4),
    .io_in_data_3_5(ffb2_io_in_data_3_5),
    .io_in_data_3_6(ffb2_io_in_data_3_6),
    .io_in_data_3_7(ffb2_io_in_data_3_7),
    .io_in_tag_0_0(ffb2_io_in_tag_0_0),
    .io_in_tag_0_1(ffb2_io_in_tag_0_1),
    .io_in_tag_0_2(ffb2_io_in_tag_0_2),
    .io_in_tag_0_3(ffb2_io_in_tag_0_3),
    .io_in_tag_0_4(ffb2_io_in_tag_0_4),
    .io_in_tag_0_5(ffb2_io_in_tag_0_5),
    .io_in_tag_0_6(ffb2_io_in_tag_0_6),
    .io_in_tag_0_7(ffb2_io_in_tag_0_7),
    .io_in_tag_1_0(ffb2_io_in_tag_1_0),
    .io_in_tag_1_1(ffb2_io_in_tag_1_1),
    .io_in_tag_1_2(ffb2_io_in_tag_1_2),
    .io_in_tag_1_3(ffb2_io_in_tag_1_3),
    .io_in_tag_1_4(ffb2_io_in_tag_1_4),
    .io_in_tag_1_5(ffb2_io_in_tag_1_5),
    .io_in_tag_1_6(ffb2_io_in_tag_1_6),
    .io_in_tag_1_7(ffb2_io_in_tag_1_7),
    .io_in_tag_2_0(ffb2_io_in_tag_2_0),
    .io_in_tag_2_1(ffb2_io_in_tag_2_1),
    .io_in_tag_2_2(ffb2_io_in_tag_2_2),
    .io_in_tag_2_3(ffb2_io_in_tag_2_3),
    .io_in_tag_2_4(ffb2_io_in_tag_2_4),
    .io_in_tag_2_5(ffb2_io_in_tag_2_5),
    .io_in_tag_2_6(ffb2_io_in_tag_2_6),
    .io_in_tag_2_7(ffb2_io_in_tag_2_7),
    .io_in_tag_3_0(ffb2_io_in_tag_3_0),
    .io_in_tag_3_1(ffb2_io_in_tag_3_1),
    .io_in_tag_3_2(ffb2_io_in_tag_3_2),
    .io_in_tag_3_3(ffb2_io_in_tag_3_3),
    .io_in_tag_3_4(ffb2_io_in_tag_3_4),
    .io_in_tag_3_5(ffb2_io_in_tag_3_5),
    .io_in_tag_3_6(ffb2_io_in_tag_3_6),
    .io_in_tag_3_7(ffb2_io_in_tag_3_7),
    .io_out_data_0_0(ffb2_io_out_data_0_0),
    .io_out_data_0_1(ffb2_io_out_data_0_1),
    .io_out_data_0_2(ffb2_io_out_data_0_2),
    .io_out_data_0_3(ffb2_io_out_data_0_3),
    .io_out_data_0_4(ffb2_io_out_data_0_4),
    .io_out_data_0_5(ffb2_io_out_data_0_5),
    .io_out_data_0_6(ffb2_io_out_data_0_6),
    .io_out_data_0_7(ffb2_io_out_data_0_7),
    .io_out_data_1_0(ffb2_io_out_data_1_0),
    .io_out_data_1_1(ffb2_io_out_data_1_1),
    .io_out_data_1_2(ffb2_io_out_data_1_2),
    .io_out_data_1_3(ffb2_io_out_data_1_3),
    .io_out_data_1_4(ffb2_io_out_data_1_4),
    .io_out_data_1_5(ffb2_io_out_data_1_5),
    .io_out_data_1_6(ffb2_io_out_data_1_6),
    .io_out_data_1_7(ffb2_io_out_data_1_7),
    .io_out_data_2_0(ffb2_io_out_data_2_0),
    .io_out_data_2_1(ffb2_io_out_data_2_1),
    .io_out_data_2_2(ffb2_io_out_data_2_2),
    .io_out_data_2_3(ffb2_io_out_data_2_3),
    .io_out_data_2_4(ffb2_io_out_data_2_4),
    .io_out_data_2_5(ffb2_io_out_data_2_5),
    .io_out_data_2_6(ffb2_io_out_data_2_6),
    .io_out_data_2_7(ffb2_io_out_data_2_7),
    .io_out_data_3_0(ffb2_io_out_data_3_0),
    .io_out_data_3_1(ffb2_io_out_data_3_1),
    .io_out_data_3_2(ffb2_io_out_data_3_2),
    .io_out_data_3_3(ffb2_io_out_data_3_3),
    .io_out_data_3_4(ffb2_io_out_data_3_4),
    .io_out_data_3_5(ffb2_io_out_data_3_5),
    .io_out_data_3_6(ffb2_io_out_data_3_6),
    .io_out_data_3_7(ffb2_io_out_data_3_7),
    .io_out_tag_0_0(ffb2_io_out_tag_0_0),
    .io_out_tag_0_1(ffb2_io_out_tag_0_1),
    .io_out_tag_0_2(ffb2_io_out_tag_0_2),
    .io_out_tag_0_3(ffb2_io_out_tag_0_3),
    .io_out_tag_0_4(ffb2_io_out_tag_0_4),
    .io_out_tag_0_5(ffb2_io_out_tag_0_5),
    .io_out_tag_0_6(ffb2_io_out_tag_0_6),
    .io_out_tag_0_7(ffb2_io_out_tag_0_7),
    .io_out_tag_1_0(ffb2_io_out_tag_1_0),
    .io_out_tag_1_1(ffb2_io_out_tag_1_1),
    .io_out_tag_1_2(ffb2_io_out_tag_1_2),
    .io_out_tag_1_3(ffb2_io_out_tag_1_3),
    .io_out_tag_1_4(ffb2_io_out_tag_1_4),
    .io_out_tag_1_5(ffb2_io_out_tag_1_5),
    .io_out_tag_1_6(ffb2_io_out_tag_1_6),
    .io_out_tag_1_7(ffb2_io_out_tag_1_7),
    .io_out_tag_2_0(ffb2_io_out_tag_2_0),
    .io_out_tag_2_1(ffb2_io_out_tag_2_1),
    .io_out_tag_2_2(ffb2_io_out_tag_2_2),
    .io_out_tag_2_3(ffb2_io_out_tag_2_3),
    .io_out_tag_2_4(ffb2_io_out_tag_2_4),
    .io_out_tag_2_5(ffb2_io_out_tag_2_5),
    .io_out_tag_2_6(ffb2_io_out_tag_2_6),
    .io_out_tag_2_7(ffb2_io_out_tag_2_7),
    .io_out_tag_3_0(ffb2_io_out_tag_3_0),
    .io_out_tag_3_1(ffb2_io_out_tag_3_1),
    .io_out_tag_3_2(ffb2_io_out_tag_3_2),
    .io_out_tag_3_3(ffb2_io_out_tag_3_3),
    .io_out_tag_3_4(ffb2_io_out_tag_3_4),
    .io_out_tag_3_5(ffb2_io_out_tag_3_5),
    .io_out_tag_3_6(ffb2_io_out_tag_3_6),
    .io_out_tag_3_7(ffb2_io_out_tag_3_7)
  );
  FF8 ffa1( // @[STA_VDBB.scala 71:20:@9792.4]
    .clock(ffa1_clock),
    .reset(ffa1_reset),
    .io_in_data_0_0(ffa1_io_in_data_0_0),
    .io_in_data_0_1(ffa1_io_in_data_0_1),
    .io_in_data_0_2(ffa1_io_in_data_0_2),
    .io_in_data_0_3(ffa1_io_in_data_0_3),
    .io_in_data_0_4(ffa1_io_in_data_0_4),
    .io_in_data_0_5(ffa1_io_in_data_0_5),
    .io_in_data_0_6(ffa1_io_in_data_0_6),
    .io_in_data_0_7(ffa1_io_in_data_0_7),
    .io_in_data_1_0(ffa1_io_in_data_1_0),
    .io_in_data_1_1(ffa1_io_in_data_1_1),
    .io_in_data_1_2(ffa1_io_in_data_1_2),
    .io_in_data_1_3(ffa1_io_in_data_1_3),
    .io_in_data_1_4(ffa1_io_in_data_1_4),
    .io_in_data_1_5(ffa1_io_in_data_1_5),
    .io_in_data_1_6(ffa1_io_in_data_1_6),
    .io_in_data_1_7(ffa1_io_in_data_1_7),
    .io_out_data_0_0(ffa1_io_out_data_0_0),
    .io_out_data_0_1(ffa1_io_out_data_0_1),
    .io_out_data_0_2(ffa1_io_out_data_0_2),
    .io_out_data_0_3(ffa1_io_out_data_0_3),
    .io_out_data_0_4(ffa1_io_out_data_0_4),
    .io_out_data_0_5(ffa1_io_out_data_0_5),
    .io_out_data_0_6(ffa1_io_out_data_0_6),
    .io_out_data_0_7(ffa1_io_out_data_0_7),
    .io_out_data_1_0(ffa1_io_out_data_1_0),
    .io_out_data_1_1(ffa1_io_out_data_1_1),
    .io_out_data_1_2(ffa1_io_out_data_1_2),
    .io_out_data_1_3(ffa1_io_out_data_1_3),
    .io_out_data_1_4(ffa1_io_out_data_1_4),
    .io_out_data_1_5(ffa1_io_out_data_1_5),
    .io_out_data_1_6(ffa1_io_out_data_1_6),
    .io_out_data_1_7(ffa1_io_out_data_1_7)
  );
  FF8 ff00( // @[STA_VDBB.scala 72:20:@9795.4]
    .clock(ff00_clock),
    .reset(ff00_reset),
    .io_in_data_0_0(ff00_io_in_data_0_0),
    .io_in_data_0_1(ff00_io_in_data_0_1),
    .io_in_data_0_2(ff00_io_in_data_0_2),
    .io_in_data_0_3(ff00_io_in_data_0_3),
    .io_in_data_0_4(ff00_io_in_data_0_4),
    .io_in_data_0_5(ff00_io_in_data_0_5),
    .io_in_data_0_6(ff00_io_in_data_0_6),
    .io_in_data_0_7(ff00_io_in_data_0_7),
    .io_in_data_1_0(ff00_io_in_data_1_0),
    .io_in_data_1_1(ff00_io_in_data_1_1),
    .io_in_data_1_2(ff00_io_in_data_1_2),
    .io_in_data_1_3(ff00_io_in_data_1_3),
    .io_in_data_1_4(ff00_io_in_data_1_4),
    .io_in_data_1_5(ff00_io_in_data_1_5),
    .io_in_data_1_6(ff00_io_in_data_1_6),
    .io_in_data_1_7(ff00_io_in_data_1_7),
    .io_out_data_0_0(ff00_io_out_data_0_0),
    .io_out_data_0_1(ff00_io_out_data_0_1),
    .io_out_data_0_2(ff00_io_out_data_0_2),
    .io_out_data_0_3(ff00_io_out_data_0_3),
    .io_out_data_0_4(ff00_io_out_data_0_4),
    .io_out_data_0_5(ff00_io_out_data_0_5),
    .io_out_data_0_6(ff00_io_out_data_0_6),
    .io_out_data_0_7(ff00_io_out_data_0_7),
    .io_out_data_1_0(ff00_io_out_data_1_0),
    .io_out_data_1_1(ff00_io_out_data_1_1),
    .io_out_data_1_2(ff00_io_out_data_1_2),
    .io_out_data_1_3(ff00_io_out_data_1_3),
    .io_out_data_1_4(ff00_io_out_data_1_4),
    .io_out_data_1_5(ff00_io_out_data_1_5),
    .io_out_data_1_6(ff00_io_out_data_1_6),
    .io_out_data_1_7(ff00_io_out_data_1_7)
  );
  FF4 ff01( // @[STA_VDBB.scala 74:20:@9798.4]
    .clock(ff01_clock),
    .reset(ff01_reset),
    .io_in_data_0_0(ff01_io_in_data_0_0),
    .io_in_data_0_1(ff01_io_in_data_0_1),
    .io_in_data_0_2(ff01_io_in_data_0_2),
    .io_in_data_0_3(ff01_io_in_data_0_3),
    .io_in_data_0_4(ff01_io_in_data_0_4),
    .io_in_data_0_5(ff01_io_in_data_0_5),
    .io_in_data_0_6(ff01_io_in_data_0_6),
    .io_in_data_0_7(ff01_io_in_data_0_7),
    .io_in_data_1_0(ff01_io_in_data_1_0),
    .io_in_data_1_1(ff01_io_in_data_1_1),
    .io_in_data_1_2(ff01_io_in_data_1_2),
    .io_in_data_1_3(ff01_io_in_data_1_3),
    .io_in_data_1_4(ff01_io_in_data_1_4),
    .io_in_data_1_5(ff01_io_in_data_1_5),
    .io_in_data_1_6(ff01_io_in_data_1_6),
    .io_in_data_1_7(ff01_io_in_data_1_7),
    .io_in_data_2_0(ff01_io_in_data_2_0),
    .io_in_data_2_1(ff01_io_in_data_2_1),
    .io_in_data_2_2(ff01_io_in_data_2_2),
    .io_in_data_2_3(ff01_io_in_data_2_3),
    .io_in_data_2_4(ff01_io_in_data_2_4),
    .io_in_data_2_5(ff01_io_in_data_2_5),
    .io_in_data_2_6(ff01_io_in_data_2_6),
    .io_in_data_2_7(ff01_io_in_data_2_7),
    .io_in_data_3_0(ff01_io_in_data_3_0),
    .io_in_data_3_1(ff01_io_in_data_3_1),
    .io_in_data_3_2(ff01_io_in_data_3_2),
    .io_in_data_3_3(ff01_io_in_data_3_3),
    .io_in_data_3_4(ff01_io_in_data_3_4),
    .io_in_data_3_5(ff01_io_in_data_3_5),
    .io_in_data_3_6(ff01_io_in_data_3_6),
    .io_in_data_3_7(ff01_io_in_data_3_7),
    .io_in_tag_0_0(ff01_io_in_tag_0_0),
    .io_in_tag_0_1(ff01_io_in_tag_0_1),
    .io_in_tag_0_2(ff01_io_in_tag_0_2),
    .io_in_tag_0_3(ff01_io_in_tag_0_3),
    .io_in_tag_0_4(ff01_io_in_tag_0_4),
    .io_in_tag_0_5(ff01_io_in_tag_0_5),
    .io_in_tag_0_6(ff01_io_in_tag_0_6),
    .io_in_tag_0_7(ff01_io_in_tag_0_7),
    .io_in_tag_1_0(ff01_io_in_tag_1_0),
    .io_in_tag_1_1(ff01_io_in_tag_1_1),
    .io_in_tag_1_2(ff01_io_in_tag_1_2),
    .io_in_tag_1_3(ff01_io_in_tag_1_3),
    .io_in_tag_1_4(ff01_io_in_tag_1_4),
    .io_in_tag_1_5(ff01_io_in_tag_1_5),
    .io_in_tag_1_6(ff01_io_in_tag_1_6),
    .io_in_tag_1_7(ff01_io_in_tag_1_7),
    .io_in_tag_2_0(ff01_io_in_tag_2_0),
    .io_in_tag_2_1(ff01_io_in_tag_2_1),
    .io_in_tag_2_2(ff01_io_in_tag_2_2),
    .io_in_tag_2_3(ff01_io_in_tag_2_3),
    .io_in_tag_2_4(ff01_io_in_tag_2_4),
    .io_in_tag_2_5(ff01_io_in_tag_2_5),
    .io_in_tag_2_6(ff01_io_in_tag_2_6),
    .io_in_tag_2_7(ff01_io_in_tag_2_7),
    .io_in_tag_3_0(ff01_io_in_tag_3_0),
    .io_in_tag_3_1(ff01_io_in_tag_3_1),
    .io_in_tag_3_2(ff01_io_in_tag_3_2),
    .io_in_tag_3_3(ff01_io_in_tag_3_3),
    .io_in_tag_3_4(ff01_io_in_tag_3_4),
    .io_in_tag_3_5(ff01_io_in_tag_3_5),
    .io_in_tag_3_6(ff01_io_in_tag_3_6),
    .io_in_tag_3_7(ff01_io_in_tag_3_7),
    .io_out_data_0_0(ff01_io_out_data_0_0),
    .io_out_data_0_1(ff01_io_out_data_0_1),
    .io_out_data_0_2(ff01_io_out_data_0_2),
    .io_out_data_0_3(ff01_io_out_data_0_3),
    .io_out_data_0_4(ff01_io_out_data_0_4),
    .io_out_data_0_5(ff01_io_out_data_0_5),
    .io_out_data_0_6(ff01_io_out_data_0_6),
    .io_out_data_0_7(ff01_io_out_data_0_7),
    .io_out_data_1_0(ff01_io_out_data_1_0),
    .io_out_data_1_1(ff01_io_out_data_1_1),
    .io_out_data_1_2(ff01_io_out_data_1_2),
    .io_out_data_1_3(ff01_io_out_data_1_3),
    .io_out_data_1_4(ff01_io_out_data_1_4),
    .io_out_data_1_5(ff01_io_out_data_1_5),
    .io_out_data_1_6(ff01_io_out_data_1_6),
    .io_out_data_1_7(ff01_io_out_data_1_7),
    .io_out_data_2_0(ff01_io_out_data_2_0),
    .io_out_data_2_1(ff01_io_out_data_2_1),
    .io_out_data_2_2(ff01_io_out_data_2_2),
    .io_out_data_2_3(ff01_io_out_data_2_3),
    .io_out_data_2_4(ff01_io_out_data_2_4),
    .io_out_data_2_5(ff01_io_out_data_2_5),
    .io_out_data_2_6(ff01_io_out_data_2_6),
    .io_out_data_2_7(ff01_io_out_data_2_7),
    .io_out_data_3_0(ff01_io_out_data_3_0),
    .io_out_data_3_1(ff01_io_out_data_3_1),
    .io_out_data_3_2(ff01_io_out_data_3_2),
    .io_out_data_3_3(ff01_io_out_data_3_3),
    .io_out_data_3_4(ff01_io_out_data_3_4),
    .io_out_data_3_5(ff01_io_out_data_3_5),
    .io_out_data_3_6(ff01_io_out_data_3_6),
    .io_out_data_3_7(ff01_io_out_data_3_7),
    .io_out_tag_0_0(ff01_io_out_tag_0_0),
    .io_out_tag_0_1(ff01_io_out_tag_0_1),
    .io_out_tag_0_2(ff01_io_out_tag_0_2),
    .io_out_tag_0_3(ff01_io_out_tag_0_3),
    .io_out_tag_0_4(ff01_io_out_tag_0_4),
    .io_out_tag_0_5(ff01_io_out_tag_0_5),
    .io_out_tag_0_6(ff01_io_out_tag_0_6),
    .io_out_tag_0_7(ff01_io_out_tag_0_7),
    .io_out_tag_1_0(ff01_io_out_tag_1_0),
    .io_out_tag_1_1(ff01_io_out_tag_1_1),
    .io_out_tag_1_2(ff01_io_out_tag_1_2),
    .io_out_tag_1_3(ff01_io_out_tag_1_3),
    .io_out_tag_1_4(ff01_io_out_tag_1_4),
    .io_out_tag_1_5(ff01_io_out_tag_1_5),
    .io_out_tag_1_6(ff01_io_out_tag_1_6),
    .io_out_tag_1_7(ff01_io_out_tag_1_7),
    .io_out_tag_2_0(ff01_io_out_tag_2_0),
    .io_out_tag_2_1(ff01_io_out_tag_2_1),
    .io_out_tag_2_2(ff01_io_out_tag_2_2),
    .io_out_tag_2_3(ff01_io_out_tag_2_3),
    .io_out_tag_2_4(ff01_io_out_tag_2_4),
    .io_out_tag_2_5(ff01_io_out_tag_2_5),
    .io_out_tag_2_6(ff01_io_out_tag_2_6),
    .io_out_tag_2_7(ff01_io_out_tag_2_7),
    .io_out_tag_3_0(ff01_io_out_tag_3_0),
    .io_out_tag_3_1(ff01_io_out_tag_3_1),
    .io_out_tag_3_2(ff01_io_out_tag_3_2),
    .io_out_tag_3_3(ff01_io_out_tag_3_3),
    .io_out_tag_3_4(ff01_io_out_tag_3_4),
    .io_out_tag_3_5(ff01_io_out_tag_3_5),
    .io_out_tag_3_6(ff01_io_out_tag_3_6),
    .io_out_tag_3_7(ff01_io_out_tag_3_7)
  );
  FF4 ff10( // @[STA_VDBB.scala 75:20:@9801.4]
    .clock(ff10_clock),
    .reset(ff10_reset),
    .io_in_data_0_0(ff10_io_in_data_0_0),
    .io_in_data_0_1(ff10_io_in_data_0_1),
    .io_in_data_0_2(ff10_io_in_data_0_2),
    .io_in_data_0_3(ff10_io_in_data_0_3),
    .io_in_data_0_4(ff10_io_in_data_0_4),
    .io_in_data_0_5(ff10_io_in_data_0_5),
    .io_in_data_0_6(ff10_io_in_data_0_6),
    .io_in_data_0_7(ff10_io_in_data_0_7),
    .io_in_data_1_0(ff10_io_in_data_1_0),
    .io_in_data_1_1(ff10_io_in_data_1_1),
    .io_in_data_1_2(ff10_io_in_data_1_2),
    .io_in_data_1_3(ff10_io_in_data_1_3),
    .io_in_data_1_4(ff10_io_in_data_1_4),
    .io_in_data_1_5(ff10_io_in_data_1_5),
    .io_in_data_1_6(ff10_io_in_data_1_6),
    .io_in_data_1_7(ff10_io_in_data_1_7),
    .io_in_data_2_0(ff10_io_in_data_2_0),
    .io_in_data_2_1(ff10_io_in_data_2_1),
    .io_in_data_2_2(ff10_io_in_data_2_2),
    .io_in_data_2_3(ff10_io_in_data_2_3),
    .io_in_data_2_4(ff10_io_in_data_2_4),
    .io_in_data_2_5(ff10_io_in_data_2_5),
    .io_in_data_2_6(ff10_io_in_data_2_6),
    .io_in_data_2_7(ff10_io_in_data_2_7),
    .io_in_data_3_0(ff10_io_in_data_3_0),
    .io_in_data_3_1(ff10_io_in_data_3_1),
    .io_in_data_3_2(ff10_io_in_data_3_2),
    .io_in_data_3_3(ff10_io_in_data_3_3),
    .io_in_data_3_4(ff10_io_in_data_3_4),
    .io_in_data_3_5(ff10_io_in_data_3_5),
    .io_in_data_3_6(ff10_io_in_data_3_6),
    .io_in_data_3_7(ff10_io_in_data_3_7),
    .io_in_tag_0_0(ff10_io_in_tag_0_0),
    .io_in_tag_0_1(ff10_io_in_tag_0_1),
    .io_in_tag_0_2(ff10_io_in_tag_0_2),
    .io_in_tag_0_3(ff10_io_in_tag_0_3),
    .io_in_tag_0_4(ff10_io_in_tag_0_4),
    .io_in_tag_0_5(ff10_io_in_tag_0_5),
    .io_in_tag_0_6(ff10_io_in_tag_0_6),
    .io_in_tag_0_7(ff10_io_in_tag_0_7),
    .io_in_tag_1_0(ff10_io_in_tag_1_0),
    .io_in_tag_1_1(ff10_io_in_tag_1_1),
    .io_in_tag_1_2(ff10_io_in_tag_1_2),
    .io_in_tag_1_3(ff10_io_in_tag_1_3),
    .io_in_tag_1_4(ff10_io_in_tag_1_4),
    .io_in_tag_1_5(ff10_io_in_tag_1_5),
    .io_in_tag_1_6(ff10_io_in_tag_1_6),
    .io_in_tag_1_7(ff10_io_in_tag_1_7),
    .io_in_tag_2_0(ff10_io_in_tag_2_0),
    .io_in_tag_2_1(ff10_io_in_tag_2_1),
    .io_in_tag_2_2(ff10_io_in_tag_2_2),
    .io_in_tag_2_3(ff10_io_in_tag_2_3),
    .io_in_tag_2_4(ff10_io_in_tag_2_4),
    .io_in_tag_2_5(ff10_io_in_tag_2_5),
    .io_in_tag_2_6(ff10_io_in_tag_2_6),
    .io_in_tag_2_7(ff10_io_in_tag_2_7),
    .io_in_tag_3_0(ff10_io_in_tag_3_0),
    .io_in_tag_3_1(ff10_io_in_tag_3_1),
    .io_in_tag_3_2(ff10_io_in_tag_3_2),
    .io_in_tag_3_3(ff10_io_in_tag_3_3),
    .io_in_tag_3_4(ff10_io_in_tag_3_4),
    .io_in_tag_3_5(ff10_io_in_tag_3_5),
    .io_in_tag_3_6(ff10_io_in_tag_3_6),
    .io_in_tag_3_7(ff10_io_in_tag_3_7),
    .io_out_data_0_0(ff10_io_out_data_0_0),
    .io_out_data_0_1(ff10_io_out_data_0_1),
    .io_out_data_0_2(ff10_io_out_data_0_2),
    .io_out_data_0_3(ff10_io_out_data_0_3),
    .io_out_data_0_4(ff10_io_out_data_0_4),
    .io_out_data_0_5(ff10_io_out_data_0_5),
    .io_out_data_0_6(ff10_io_out_data_0_6),
    .io_out_data_0_7(ff10_io_out_data_0_7),
    .io_out_data_1_0(ff10_io_out_data_1_0),
    .io_out_data_1_1(ff10_io_out_data_1_1),
    .io_out_data_1_2(ff10_io_out_data_1_2),
    .io_out_data_1_3(ff10_io_out_data_1_3),
    .io_out_data_1_4(ff10_io_out_data_1_4),
    .io_out_data_1_5(ff10_io_out_data_1_5),
    .io_out_data_1_6(ff10_io_out_data_1_6),
    .io_out_data_1_7(ff10_io_out_data_1_7),
    .io_out_data_2_0(ff10_io_out_data_2_0),
    .io_out_data_2_1(ff10_io_out_data_2_1),
    .io_out_data_2_2(ff10_io_out_data_2_2),
    .io_out_data_2_3(ff10_io_out_data_2_3),
    .io_out_data_2_4(ff10_io_out_data_2_4),
    .io_out_data_2_5(ff10_io_out_data_2_5),
    .io_out_data_2_6(ff10_io_out_data_2_6),
    .io_out_data_2_7(ff10_io_out_data_2_7),
    .io_out_data_3_0(ff10_io_out_data_3_0),
    .io_out_data_3_1(ff10_io_out_data_3_1),
    .io_out_data_3_2(ff10_io_out_data_3_2),
    .io_out_data_3_3(ff10_io_out_data_3_3),
    .io_out_data_3_4(ff10_io_out_data_3_4),
    .io_out_data_3_5(ff10_io_out_data_3_5),
    .io_out_data_3_6(ff10_io_out_data_3_6),
    .io_out_data_3_7(ff10_io_out_data_3_7),
    .io_out_tag_0_0(ff10_io_out_tag_0_0),
    .io_out_tag_0_1(ff10_io_out_tag_0_1),
    .io_out_tag_0_2(ff10_io_out_tag_0_2),
    .io_out_tag_0_3(ff10_io_out_tag_0_3),
    .io_out_tag_0_4(ff10_io_out_tag_0_4),
    .io_out_tag_0_5(ff10_io_out_tag_0_5),
    .io_out_tag_0_6(ff10_io_out_tag_0_6),
    .io_out_tag_0_7(ff10_io_out_tag_0_7),
    .io_out_tag_1_0(ff10_io_out_tag_1_0),
    .io_out_tag_1_1(ff10_io_out_tag_1_1),
    .io_out_tag_1_2(ff10_io_out_tag_1_2),
    .io_out_tag_1_3(ff10_io_out_tag_1_3),
    .io_out_tag_1_4(ff10_io_out_tag_1_4),
    .io_out_tag_1_5(ff10_io_out_tag_1_5),
    .io_out_tag_1_6(ff10_io_out_tag_1_6),
    .io_out_tag_1_7(ff10_io_out_tag_1_7),
    .io_out_tag_2_0(ff10_io_out_tag_2_0),
    .io_out_tag_2_1(ff10_io_out_tag_2_1),
    .io_out_tag_2_2(ff10_io_out_tag_2_2),
    .io_out_tag_2_3(ff10_io_out_tag_2_3),
    .io_out_tag_2_4(ff10_io_out_tag_2_4),
    .io_out_tag_2_5(ff10_io_out_tag_2_5),
    .io_out_tag_2_6(ff10_io_out_tag_2_6),
    .io_out_tag_2_7(ff10_io_out_tag_2_7),
    .io_out_tag_3_0(ff10_io_out_tag_3_0),
    .io_out_tag_3_1(ff10_io_out_tag_3_1),
    .io_out_tag_3_2(ff10_io_out_tag_3_2),
    .io_out_tag_3_3(ff10_io_out_tag_3_3),
    .io_out_tag_3_4(ff10_io_out_tag_3_4),
    .io_out_tag_3_5(ff10_io_out_tag_3_5),
    .io_out_tag_3_6(ff10_io_out_tag_3_6),
    .io_out_tag_3_7(ff10_io_out_tag_3_7)
  );
  FF8 ffa2( // @[STA_VDBB.scala 77:20:@9804.4]
    .clock(ffa2_clock),
    .reset(ffa2_reset),
    .io_in_data_0_0(ffa2_io_in_data_0_0),
    .io_in_data_0_1(ffa2_io_in_data_0_1),
    .io_in_data_0_2(ffa2_io_in_data_0_2),
    .io_in_data_0_3(ffa2_io_in_data_0_3),
    .io_in_data_0_4(ffa2_io_in_data_0_4),
    .io_in_data_0_5(ffa2_io_in_data_0_5),
    .io_in_data_0_6(ffa2_io_in_data_0_6),
    .io_in_data_0_7(ffa2_io_in_data_0_7),
    .io_in_data_1_0(ffa2_io_in_data_1_0),
    .io_in_data_1_1(ffa2_io_in_data_1_1),
    .io_in_data_1_2(ffa2_io_in_data_1_2),
    .io_in_data_1_3(ffa2_io_in_data_1_3),
    .io_in_data_1_4(ffa2_io_in_data_1_4),
    .io_in_data_1_5(ffa2_io_in_data_1_5),
    .io_in_data_1_6(ffa2_io_in_data_1_6),
    .io_in_data_1_7(ffa2_io_in_data_1_7),
    .io_out_data_0_0(ffa2_io_out_data_0_0),
    .io_out_data_0_1(ffa2_io_out_data_0_1),
    .io_out_data_0_2(ffa2_io_out_data_0_2),
    .io_out_data_0_3(ffa2_io_out_data_0_3),
    .io_out_data_0_4(ffa2_io_out_data_0_4),
    .io_out_data_0_5(ffa2_io_out_data_0_5),
    .io_out_data_0_6(ffa2_io_out_data_0_6),
    .io_out_data_0_7(ffa2_io_out_data_0_7),
    .io_out_data_1_0(ffa2_io_out_data_1_0),
    .io_out_data_1_1(ffa2_io_out_data_1_1),
    .io_out_data_1_2(ffa2_io_out_data_1_2),
    .io_out_data_1_3(ffa2_io_out_data_1_3),
    .io_out_data_1_4(ffa2_io_out_data_1_4),
    .io_out_data_1_5(ffa2_io_out_data_1_5),
    .io_out_data_1_6(ffa2_io_out_data_1_6),
    .io_out_data_1_7(ffa2_io_out_data_1_7)
  );
  FF8 ff11( // @[STA_VDBB.scala 78:20:@9807.4]
    .clock(ff11_clock),
    .reset(ff11_reset),
    .io_in_data_0_0(ff11_io_in_data_0_0),
    .io_in_data_0_1(ff11_io_in_data_0_1),
    .io_in_data_0_2(ff11_io_in_data_0_2),
    .io_in_data_0_3(ff11_io_in_data_0_3),
    .io_in_data_0_4(ff11_io_in_data_0_4),
    .io_in_data_0_5(ff11_io_in_data_0_5),
    .io_in_data_0_6(ff11_io_in_data_0_6),
    .io_in_data_0_7(ff11_io_in_data_0_7),
    .io_in_data_1_0(ff11_io_in_data_1_0),
    .io_in_data_1_1(ff11_io_in_data_1_1),
    .io_in_data_1_2(ff11_io_in_data_1_2),
    .io_in_data_1_3(ff11_io_in_data_1_3),
    .io_in_data_1_4(ff11_io_in_data_1_4),
    .io_in_data_1_5(ff11_io_in_data_1_5),
    .io_in_data_1_6(ff11_io_in_data_1_6),
    .io_in_data_1_7(ff11_io_in_data_1_7),
    .io_out_data_0_0(ff11_io_out_data_0_0),
    .io_out_data_0_1(ff11_io_out_data_0_1),
    .io_out_data_0_2(ff11_io_out_data_0_2),
    .io_out_data_0_3(ff11_io_out_data_0_3),
    .io_out_data_0_4(ff11_io_out_data_0_4),
    .io_out_data_0_5(ff11_io_out_data_0_5),
    .io_out_data_0_6(ff11_io_out_data_0_6),
    .io_out_data_0_7(ff11_io_out_data_0_7),
    .io_out_data_1_0(ff11_io_out_data_1_0),
    .io_out_data_1_1(ff11_io_out_data_1_1),
    .io_out_data_1_2(ff11_io_out_data_1_2),
    .io_out_data_1_3(ff11_io_out_data_1_3),
    .io_out_data_1_4(ff11_io_out_data_1_4),
    .io_out_data_1_5(ff11_io_out_data_1_5),
    .io_out_data_1_6(ff11_io_out_data_1_6),
    .io_out_data_1_7(ff11_io_out_data_1_7)
  );
  assign S8DP1s_0_0_result = S8DP1_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8879.4]
  assign S8DP1s_0_1_result = S8DP1_1_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8905.4]
  assign S8DP1s_0_2_result = S8DP1_2_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8931.4]
  assign S8DP1s_0_3_result = S8DP1_3_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8957.4]
  assign S8DP1s_0_4_result = S8DP1_4_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@8983.4]
  assign S8DP1s_0_5_result = S8DP1_5_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9009.4]
  assign S8DP1s_0_6_result = S8DP1_6_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9035.4]
  assign S8DP1s_0_7_result = S8DP1_7_io_result; // @[STA_VDBB.scala 55:21:@8878.4 STA_VDBB.scala 55:21:@9061.4]
  assign S8DP1s_1_0_result = S8DP1_8_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9112.4]
  assign S8DP1s_1_1_result = S8DP1_9_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9138.4]
  assign S8DP1s_1_2_result = S8DP1_10_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9164.4]
  assign S8DP1s_1_3_result = S8DP1_11_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9190.4]
  assign S8DP1s_1_4_result = S8DP1_12_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9216.4]
  assign S8DP1s_1_5_result = S8DP1_13_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9242.4]
  assign S8DP1s_1_6_result = S8DP1_14_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9268.4]
  assign S8DP1s_1_7_result = S8DP1_15_io_result; // @[STA_VDBB.scala 56:21:@9111.4 STA_VDBB.scala 56:21:@9294.4]
  assign S8DP1s_2_0_result = S8DP1_16_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9345.4]
  assign S8DP1s_2_1_result = S8DP1_17_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9371.4]
  assign S8DP1s_2_2_result = S8DP1_18_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9397.4]
  assign S8DP1s_2_3_result = S8DP1_19_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9423.4]
  assign S8DP1s_2_4_result = S8DP1_20_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9449.4]
  assign S8DP1s_2_5_result = S8DP1_21_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9475.4]
  assign S8DP1s_2_6_result = S8DP1_22_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9501.4]
  assign S8DP1s_2_7_result = S8DP1_23_io_result; // @[STA_VDBB.scala 57:21:@9344.4 STA_VDBB.scala 57:21:@9527.4]
  assign S8DP1s_3_0_result = S8DP1_24_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9578.4]
  assign S8DP1s_3_1_result = S8DP1_25_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9604.4]
  assign S8DP1s_3_2_result = S8DP1_26_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9630.4]
  assign S8DP1s_3_3_result = S8DP1_27_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9656.4]
  assign S8DP1s_3_4_result = S8DP1_28_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9682.4]
  assign S8DP1s_3_5_result = S8DP1_29_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9708.4]
  assign S8DP1s_3_6_result = S8DP1_30_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9734.4]
  assign S8DP1s_3_7_result = S8DP1_31_io_result; // @[STA_VDBB.scala 58:21:@9577.4 STA_VDBB.scala 58:21:@9760.4]
  assign io_out_C_0_0 = out_result_0_0; // @[STA_VDBB.scala 354:12:@27842.4]
  assign io_out_C_0_1 = out_result_0_1; // @[STA_VDBB.scala 354:12:@27843.4]
  assign io_out_C_0_2 = out_result_0_2; // @[STA_VDBB.scala 354:12:@27844.4]
  assign io_out_C_0_3 = out_result_0_3; // @[STA_VDBB.scala 354:12:@27845.4]
  assign io_out_C_0_4 = out_result_0_4; // @[STA_VDBB.scala 354:12:@27846.4]
  assign io_out_C_0_5 = out_result_0_5; // @[STA_VDBB.scala 354:12:@27847.4]
  assign io_out_C_0_6 = out_result_0_6; // @[STA_VDBB.scala 354:12:@27848.4]
  assign io_out_C_0_7 = out_result_0_7; // @[STA_VDBB.scala 354:12:@27849.4]
  assign io_out_C_1_0 = out_result_1_0; // @[STA_VDBB.scala 354:12:@27850.4]
  assign io_out_C_1_1 = out_result_1_1; // @[STA_VDBB.scala 354:12:@27851.4]
  assign io_out_C_1_2 = out_result_1_2; // @[STA_VDBB.scala 354:12:@27852.4]
  assign io_out_C_1_3 = out_result_1_3; // @[STA_VDBB.scala 354:12:@27853.4]
  assign io_out_C_1_4 = out_result_1_4; // @[STA_VDBB.scala 354:12:@27854.4]
  assign io_out_C_1_5 = out_result_1_5; // @[STA_VDBB.scala 354:12:@27855.4]
  assign io_out_C_1_6 = out_result_1_6; // @[STA_VDBB.scala 354:12:@27856.4]
  assign io_out_C_1_7 = out_result_1_7; // @[STA_VDBB.scala 354:12:@27857.4]
  assign io_out_C_2_0 = out_result_2_0; // @[STA_VDBB.scala 354:12:@27858.4]
  assign io_out_C_2_1 = out_result_2_1; // @[STA_VDBB.scala 354:12:@27859.4]
  assign io_out_C_2_2 = out_result_2_2; // @[STA_VDBB.scala 354:12:@27860.4]
  assign io_out_C_2_3 = out_result_2_3; // @[STA_VDBB.scala 354:12:@27861.4]
  assign io_out_C_2_4 = out_result_2_4; // @[STA_VDBB.scala 354:12:@27862.4]
  assign io_out_C_2_5 = out_result_2_5; // @[STA_VDBB.scala 354:12:@27863.4]
  assign io_out_C_2_6 = out_result_2_6; // @[STA_VDBB.scala 354:12:@27864.4]
  assign io_out_C_2_7 = out_result_2_7; // @[STA_VDBB.scala 354:12:@27865.4]
  assign io_out_C_3_0 = out_result_3_0; // @[STA_VDBB.scala 354:12:@27866.4]
  assign io_out_C_3_1 = out_result_3_1; // @[STA_VDBB.scala 354:12:@27867.4]
  assign io_out_C_3_2 = out_result_3_2; // @[STA_VDBB.scala 354:12:@27868.4]
  assign io_out_C_3_3 = out_result_3_3; // @[STA_VDBB.scala 354:12:@27869.4]
  assign io_out_C_3_4 = out_result_3_4; // @[STA_VDBB.scala 354:12:@27870.4]
  assign io_out_C_3_5 = out_result_3_5; // @[STA_VDBB.scala 354:12:@27871.4]
  assign io_out_C_3_6 = out_result_3_6; // @[STA_VDBB.scala 354:12:@27872.4]
  assign io_out_C_3_7 = out_result_3_7; // @[STA_VDBB.scala 354:12:@27873.4]
  assign tag_clock = clock; // @[:@8693.4]
  assign tag_reset = reset; // @[:@8694.4]
  assign tag_1_clock = clock; // @[:@8696.4]
  assign tag_1_reset = reset; // @[:@8697.4]
  assign tag_2_clock = clock; // @[:@8699.4]
  assign tag_2_reset = reset; // @[:@8700.4]
  assign tag_3_clock = clock; // @[:@8702.4]
  assign tag_3_reset = reset; // @[:@8703.4]
  assign MUX8_io_int_in_0 = ff10_io_out_data_0_0; // @[STA_VDBB.scala 52:17:@8795.4]
  assign MUX8_io_int_in_1 = ff10_io_out_data_0_1; // @[STA_VDBB.scala 52:17:@8796.4]
  assign MUX8_io_int_in_2 = ff10_io_out_data_0_2; // @[STA_VDBB.scala 52:17:@8797.4]
  assign MUX8_io_int_in_3 = ff10_io_out_data_0_3; // @[STA_VDBB.scala 52:17:@8798.4]
  assign MUX8_io_int_in_4 = ff10_io_out_data_0_4; // @[STA_VDBB.scala 52:17:@8799.4]
  assign MUX8_io_int_in_5 = ff10_io_out_data_0_5; // @[STA_VDBB.scala 52:17:@8800.4]
  assign MUX8_io_int_in_6 = ff10_io_out_data_0_6; // @[STA_VDBB.scala 52:17:@8801.4]
  assign MUX8_io_int_in_7 = ff10_io_out_data_0_7; // @[STA_VDBB.scala 52:17:@8802.4]
  assign MUX8_io_tag_0 = ff10_io_out_tag_0_0; // @[STA_VDBB.scala 52:17:@8787.4]
  assign MUX8_io_tag_1 = ff10_io_out_tag_0_1; // @[STA_VDBB.scala 52:17:@8788.4]
  assign MUX8_io_tag_2 = ff10_io_out_tag_0_2; // @[STA_VDBB.scala 52:17:@8789.4]
  assign MUX8_io_tag_3 = ff10_io_out_tag_0_3; // @[STA_VDBB.scala 52:17:@8790.4]
  assign MUX8_io_tag_4 = ff10_io_out_tag_0_4; // @[STA_VDBB.scala 52:17:@8791.4]
  assign MUX8_io_tag_5 = ff10_io_out_tag_0_5; // @[STA_VDBB.scala 52:17:@8792.4]
  assign MUX8_io_tag_6 = ff10_io_out_tag_0_6; // @[STA_VDBB.scala 52:17:@8793.4]
  assign MUX8_io_tag_7 = ff10_io_out_tag_0_7; // @[STA_VDBB.scala 52:17:@8794.4]
  assign MUX8_1_io_int_in_0 = ff10_io_out_data_1_0; // @[STA_VDBB.scala 52:17:@8812.4]
  assign MUX8_1_io_int_in_1 = ff10_io_out_data_1_1; // @[STA_VDBB.scala 52:17:@8813.4]
  assign MUX8_1_io_int_in_2 = ff10_io_out_data_1_2; // @[STA_VDBB.scala 52:17:@8814.4]
  assign MUX8_1_io_int_in_3 = ff10_io_out_data_1_3; // @[STA_VDBB.scala 52:17:@8815.4]
  assign MUX8_1_io_int_in_4 = ff10_io_out_data_1_4; // @[STA_VDBB.scala 52:17:@8816.4]
  assign MUX8_1_io_int_in_5 = ff10_io_out_data_1_5; // @[STA_VDBB.scala 52:17:@8817.4]
  assign MUX8_1_io_int_in_6 = ff10_io_out_data_1_6; // @[STA_VDBB.scala 52:17:@8818.4]
  assign MUX8_1_io_int_in_7 = ff10_io_out_data_1_7; // @[STA_VDBB.scala 52:17:@8819.4]
  assign MUX8_1_io_tag_0 = ff10_io_out_tag_1_0; // @[STA_VDBB.scala 52:17:@8804.4]
  assign MUX8_1_io_tag_1 = ff10_io_out_tag_1_1; // @[STA_VDBB.scala 52:17:@8805.4]
  assign MUX8_1_io_tag_2 = ff10_io_out_tag_1_2; // @[STA_VDBB.scala 52:17:@8806.4]
  assign MUX8_1_io_tag_3 = ff10_io_out_tag_1_3; // @[STA_VDBB.scala 52:17:@8807.4]
  assign MUX8_1_io_tag_4 = ff10_io_out_tag_1_4; // @[STA_VDBB.scala 52:17:@8808.4]
  assign MUX8_1_io_tag_5 = ff10_io_out_tag_1_5; // @[STA_VDBB.scala 52:17:@8809.4]
  assign MUX8_1_io_tag_6 = ff10_io_out_tag_1_6; // @[STA_VDBB.scala 52:17:@8810.4]
  assign MUX8_1_io_tag_7 = ff10_io_out_tag_1_7; // @[STA_VDBB.scala 52:17:@8811.4]
  assign MUX8_2_io_int_in_0 = ff10_io_out_data_2_0; // @[STA_VDBB.scala 52:17:@8829.4]
  assign MUX8_2_io_int_in_1 = ff10_io_out_data_2_1; // @[STA_VDBB.scala 52:17:@8830.4]
  assign MUX8_2_io_int_in_2 = ff10_io_out_data_2_2; // @[STA_VDBB.scala 52:17:@8831.4]
  assign MUX8_2_io_int_in_3 = ff10_io_out_data_2_3; // @[STA_VDBB.scala 52:17:@8832.4]
  assign MUX8_2_io_int_in_4 = ff10_io_out_data_2_4; // @[STA_VDBB.scala 52:17:@8833.4]
  assign MUX8_2_io_int_in_5 = ff10_io_out_data_2_5; // @[STA_VDBB.scala 52:17:@8834.4]
  assign MUX8_2_io_int_in_6 = ff10_io_out_data_2_6; // @[STA_VDBB.scala 52:17:@8835.4]
  assign MUX8_2_io_int_in_7 = ff10_io_out_data_2_7; // @[STA_VDBB.scala 52:17:@8836.4]
  assign MUX8_2_io_tag_0 = ff10_io_out_tag_2_0; // @[STA_VDBB.scala 52:17:@8821.4]
  assign MUX8_2_io_tag_1 = ff10_io_out_tag_2_1; // @[STA_VDBB.scala 52:17:@8822.4]
  assign MUX8_2_io_tag_2 = ff10_io_out_tag_2_2; // @[STA_VDBB.scala 52:17:@8823.4]
  assign MUX8_2_io_tag_3 = ff10_io_out_tag_2_3; // @[STA_VDBB.scala 52:17:@8824.4]
  assign MUX8_2_io_tag_4 = ff10_io_out_tag_2_4; // @[STA_VDBB.scala 52:17:@8825.4]
  assign MUX8_2_io_tag_5 = ff10_io_out_tag_2_5; // @[STA_VDBB.scala 52:17:@8826.4]
  assign MUX8_2_io_tag_6 = ff10_io_out_tag_2_6; // @[STA_VDBB.scala 52:17:@8827.4]
  assign MUX8_2_io_tag_7 = ff10_io_out_tag_2_7; // @[STA_VDBB.scala 52:17:@8828.4]
  assign MUX8_3_io_int_in_0 = ff10_io_out_data_3_0; // @[STA_VDBB.scala 52:17:@8846.4]
  assign MUX8_3_io_int_in_1 = ff10_io_out_data_3_1; // @[STA_VDBB.scala 52:17:@8847.4]
  assign MUX8_3_io_int_in_2 = ff10_io_out_data_3_2; // @[STA_VDBB.scala 52:17:@8848.4]
  assign MUX8_3_io_int_in_3 = ff10_io_out_data_3_3; // @[STA_VDBB.scala 52:17:@8849.4]
  assign MUX8_3_io_int_in_4 = ff10_io_out_data_3_4; // @[STA_VDBB.scala 52:17:@8850.4]
  assign MUX8_3_io_int_in_5 = ff10_io_out_data_3_5; // @[STA_VDBB.scala 52:17:@8851.4]
  assign MUX8_3_io_int_in_6 = ff10_io_out_data_3_6; // @[STA_VDBB.scala 52:17:@8852.4]
  assign MUX8_3_io_int_in_7 = ff10_io_out_data_3_7; // @[STA_VDBB.scala 52:17:@8853.4]
  assign MUX8_3_io_tag_0 = ff10_io_out_tag_3_0; // @[STA_VDBB.scala 52:17:@8838.4]
  assign MUX8_3_io_tag_1 = ff10_io_out_tag_3_1; // @[STA_VDBB.scala 52:17:@8839.4]
  assign MUX8_3_io_tag_2 = ff10_io_out_tag_3_2; // @[STA_VDBB.scala 52:17:@8840.4]
  assign MUX8_3_io_tag_3 = ff10_io_out_tag_3_3; // @[STA_VDBB.scala 52:17:@8841.4]
  assign MUX8_3_io_tag_4 = ff10_io_out_tag_3_4; // @[STA_VDBB.scala 52:17:@8842.4]
  assign MUX8_3_io_tag_5 = ff10_io_out_tag_3_5; // @[STA_VDBB.scala 52:17:@8843.4]
  assign MUX8_3_io_tag_6 = ff10_io_out_tag_3_6; // @[STA_VDBB.scala 52:17:@8844.4]
  assign MUX8_3_io_tag_7 = ff10_io_out_tag_3_7; // @[STA_VDBB.scala 52:17:@8845.4]
  assign S8DP1_clock = clock; // @[:@8855.4]
  assign S8DP1_reset = reset; // @[:@8856.4]
  assign S8DP1_io_int_in_A_0 = ffa1_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@8897.4]
  assign S8DP1_io_int_in_A_1 = ffa1_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@8898.4]
  assign S8DP1_io_int_in_A_2 = ffa1_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@8899.4]
  assign S8DP1_io_int_in_A_3 = ffa1_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@8900.4]
  assign S8DP1_io_int_in_A_4 = ffa1_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@8901.4]
  assign S8DP1_io_int_in_A_5 = ffa1_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@8902.4]
  assign S8DP1_io_int_in_A_6 = ffa1_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@8903.4]
  assign S8DP1_io_int_in_A_7 = ffa1_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@8904.4]
  assign S8DP1_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 55:21:@8896.4]
  assign S8DP1_io_tag_0 = ffb1_io_out_tag_0_0; // @[STA_VDBB.scala 55:21:@8888.4]
  assign S8DP1_io_tag_1 = ffb1_io_out_tag_0_1; // @[STA_VDBB.scala 55:21:@8889.4]
  assign S8DP1_io_tag_2 = ffb1_io_out_tag_0_2; // @[STA_VDBB.scala 55:21:@8890.4]
  assign S8DP1_io_tag_3 = ffb1_io_out_tag_0_3; // @[STA_VDBB.scala 55:21:@8891.4]
  assign S8DP1_io_tag_4 = ffb1_io_out_tag_0_4; // @[STA_VDBB.scala 55:21:@8892.4]
  assign S8DP1_io_tag_5 = ffb1_io_out_tag_0_5; // @[STA_VDBB.scala 55:21:@8893.4]
  assign S8DP1_io_tag_6 = ffb1_io_out_tag_0_6; // @[STA_VDBB.scala 55:21:@8894.4]
  assign S8DP1_io_tag_7 = ffb1_io_out_tag_0_7; // @[STA_VDBB.scala 55:21:@8895.4]
  assign S8DP1_1_clock = clock; // @[:@8858.4]
  assign S8DP1_1_reset = reset; // @[:@8859.4]
  assign S8DP1_1_io_int_in_A_0 = ffa1_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@8923.4]
  assign S8DP1_1_io_int_in_A_1 = ffa1_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@8924.4]
  assign S8DP1_1_io_int_in_A_2 = ffa1_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@8925.4]
  assign S8DP1_1_io_int_in_A_3 = ffa1_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@8926.4]
  assign S8DP1_1_io_int_in_A_4 = ffa1_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@8927.4]
  assign S8DP1_1_io_int_in_A_5 = ffa1_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@8928.4]
  assign S8DP1_1_io_int_in_A_6 = ffa1_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@8929.4]
  assign S8DP1_1_io_int_in_A_7 = ffa1_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@8930.4]
  assign S8DP1_1_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 55:21:@8922.4]
  assign S8DP1_1_io_tag_0 = ffb1_io_out_tag_1_0; // @[STA_VDBB.scala 55:21:@8914.4]
  assign S8DP1_1_io_tag_1 = ffb1_io_out_tag_1_1; // @[STA_VDBB.scala 55:21:@8915.4]
  assign S8DP1_1_io_tag_2 = ffb1_io_out_tag_1_2; // @[STA_VDBB.scala 55:21:@8916.4]
  assign S8DP1_1_io_tag_3 = ffb1_io_out_tag_1_3; // @[STA_VDBB.scala 55:21:@8917.4]
  assign S8DP1_1_io_tag_4 = ffb1_io_out_tag_1_4; // @[STA_VDBB.scala 55:21:@8918.4]
  assign S8DP1_1_io_tag_5 = ffb1_io_out_tag_1_5; // @[STA_VDBB.scala 55:21:@8919.4]
  assign S8DP1_1_io_tag_6 = ffb1_io_out_tag_1_6; // @[STA_VDBB.scala 55:21:@8920.4]
  assign S8DP1_1_io_tag_7 = ffb1_io_out_tag_1_7; // @[STA_VDBB.scala 55:21:@8921.4]
  assign S8DP1_2_clock = clock; // @[:@8861.4]
  assign S8DP1_2_reset = reset; // @[:@8862.4]
  assign S8DP1_2_io_int_in_A_0 = ffa1_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@8949.4]
  assign S8DP1_2_io_int_in_A_1 = ffa1_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@8950.4]
  assign S8DP1_2_io_int_in_A_2 = ffa1_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@8951.4]
  assign S8DP1_2_io_int_in_A_3 = ffa1_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@8952.4]
  assign S8DP1_2_io_int_in_A_4 = ffa1_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@8953.4]
  assign S8DP1_2_io_int_in_A_5 = ffa1_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@8954.4]
  assign S8DP1_2_io_int_in_A_6 = ffa1_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@8955.4]
  assign S8DP1_2_io_int_in_A_7 = ffa1_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@8956.4]
  assign S8DP1_2_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 55:21:@8948.4]
  assign S8DP1_2_io_tag_0 = ffb1_io_out_tag_2_0; // @[STA_VDBB.scala 55:21:@8940.4]
  assign S8DP1_2_io_tag_1 = ffb1_io_out_tag_2_1; // @[STA_VDBB.scala 55:21:@8941.4]
  assign S8DP1_2_io_tag_2 = ffb1_io_out_tag_2_2; // @[STA_VDBB.scala 55:21:@8942.4]
  assign S8DP1_2_io_tag_3 = ffb1_io_out_tag_2_3; // @[STA_VDBB.scala 55:21:@8943.4]
  assign S8DP1_2_io_tag_4 = ffb1_io_out_tag_2_4; // @[STA_VDBB.scala 55:21:@8944.4]
  assign S8DP1_2_io_tag_5 = ffb1_io_out_tag_2_5; // @[STA_VDBB.scala 55:21:@8945.4]
  assign S8DP1_2_io_tag_6 = ffb1_io_out_tag_2_6; // @[STA_VDBB.scala 55:21:@8946.4]
  assign S8DP1_2_io_tag_7 = ffb1_io_out_tag_2_7; // @[STA_VDBB.scala 55:21:@8947.4]
  assign S8DP1_3_clock = clock; // @[:@8864.4]
  assign S8DP1_3_reset = reset; // @[:@8865.4]
  assign S8DP1_3_io_int_in_A_0 = ffa1_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@8975.4]
  assign S8DP1_3_io_int_in_A_1 = ffa1_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@8976.4]
  assign S8DP1_3_io_int_in_A_2 = ffa1_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@8977.4]
  assign S8DP1_3_io_int_in_A_3 = ffa1_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@8978.4]
  assign S8DP1_3_io_int_in_A_4 = ffa1_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@8979.4]
  assign S8DP1_3_io_int_in_A_5 = ffa1_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@8980.4]
  assign S8DP1_3_io_int_in_A_6 = ffa1_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@8981.4]
  assign S8DP1_3_io_int_in_A_7 = ffa1_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@8982.4]
  assign S8DP1_3_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 55:21:@8974.4]
  assign S8DP1_3_io_tag_0 = ffb1_io_out_tag_3_0; // @[STA_VDBB.scala 55:21:@8966.4]
  assign S8DP1_3_io_tag_1 = ffb1_io_out_tag_3_1; // @[STA_VDBB.scala 55:21:@8967.4]
  assign S8DP1_3_io_tag_2 = ffb1_io_out_tag_3_2; // @[STA_VDBB.scala 55:21:@8968.4]
  assign S8DP1_3_io_tag_3 = ffb1_io_out_tag_3_3; // @[STA_VDBB.scala 55:21:@8969.4]
  assign S8DP1_3_io_tag_4 = ffb1_io_out_tag_3_4; // @[STA_VDBB.scala 55:21:@8970.4]
  assign S8DP1_3_io_tag_5 = ffb1_io_out_tag_3_5; // @[STA_VDBB.scala 55:21:@8971.4]
  assign S8DP1_3_io_tag_6 = ffb1_io_out_tag_3_6; // @[STA_VDBB.scala 55:21:@8972.4]
  assign S8DP1_3_io_tag_7 = ffb1_io_out_tag_3_7; // @[STA_VDBB.scala 55:21:@8973.4]
  assign S8DP1_4_clock = clock; // @[:@8867.4]
  assign S8DP1_4_reset = reset; // @[:@8868.4]
  assign S8DP1_4_io_int_in_A_0 = ff00_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@9001.4]
  assign S8DP1_4_io_int_in_A_1 = ff00_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@9002.4]
  assign S8DP1_4_io_int_in_A_2 = ff00_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@9003.4]
  assign S8DP1_4_io_int_in_A_3 = ff00_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@9004.4]
  assign S8DP1_4_io_int_in_A_4 = ff00_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@9005.4]
  assign S8DP1_4_io_int_in_A_5 = ff00_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@9006.4]
  assign S8DP1_4_io_int_in_A_6 = ff00_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@9007.4]
  assign S8DP1_4_io_int_in_A_7 = ff00_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@9008.4]
  assign S8DP1_4_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 55:21:@9000.4]
  assign S8DP1_4_io_tag_0 = ffb2_io_out_tag_0_0; // @[STA_VDBB.scala 55:21:@8992.4]
  assign S8DP1_4_io_tag_1 = ffb2_io_out_tag_0_1; // @[STA_VDBB.scala 55:21:@8993.4]
  assign S8DP1_4_io_tag_2 = ffb2_io_out_tag_0_2; // @[STA_VDBB.scala 55:21:@8994.4]
  assign S8DP1_4_io_tag_3 = ffb2_io_out_tag_0_3; // @[STA_VDBB.scala 55:21:@8995.4]
  assign S8DP1_4_io_tag_4 = ffb2_io_out_tag_0_4; // @[STA_VDBB.scala 55:21:@8996.4]
  assign S8DP1_4_io_tag_5 = ffb2_io_out_tag_0_5; // @[STA_VDBB.scala 55:21:@8997.4]
  assign S8DP1_4_io_tag_6 = ffb2_io_out_tag_0_6; // @[STA_VDBB.scala 55:21:@8998.4]
  assign S8DP1_4_io_tag_7 = ffb2_io_out_tag_0_7; // @[STA_VDBB.scala 55:21:@8999.4]
  assign S8DP1_5_clock = clock; // @[:@8870.4]
  assign S8DP1_5_reset = reset; // @[:@8871.4]
  assign S8DP1_5_io_int_in_A_0 = ff00_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@9027.4]
  assign S8DP1_5_io_int_in_A_1 = ff00_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@9028.4]
  assign S8DP1_5_io_int_in_A_2 = ff00_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@9029.4]
  assign S8DP1_5_io_int_in_A_3 = ff00_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@9030.4]
  assign S8DP1_5_io_int_in_A_4 = ff00_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@9031.4]
  assign S8DP1_5_io_int_in_A_5 = ff00_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@9032.4]
  assign S8DP1_5_io_int_in_A_6 = ff00_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@9033.4]
  assign S8DP1_5_io_int_in_A_7 = ff00_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@9034.4]
  assign S8DP1_5_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 55:21:@9026.4]
  assign S8DP1_5_io_tag_0 = ffb2_io_out_tag_1_0; // @[STA_VDBB.scala 55:21:@9018.4]
  assign S8DP1_5_io_tag_1 = ffb2_io_out_tag_1_1; // @[STA_VDBB.scala 55:21:@9019.4]
  assign S8DP1_5_io_tag_2 = ffb2_io_out_tag_1_2; // @[STA_VDBB.scala 55:21:@9020.4]
  assign S8DP1_5_io_tag_3 = ffb2_io_out_tag_1_3; // @[STA_VDBB.scala 55:21:@9021.4]
  assign S8DP1_5_io_tag_4 = ffb2_io_out_tag_1_4; // @[STA_VDBB.scala 55:21:@9022.4]
  assign S8DP1_5_io_tag_5 = ffb2_io_out_tag_1_5; // @[STA_VDBB.scala 55:21:@9023.4]
  assign S8DP1_5_io_tag_6 = ffb2_io_out_tag_1_6; // @[STA_VDBB.scala 55:21:@9024.4]
  assign S8DP1_5_io_tag_7 = ffb2_io_out_tag_1_7; // @[STA_VDBB.scala 55:21:@9025.4]
  assign S8DP1_6_clock = clock; // @[:@8873.4]
  assign S8DP1_6_reset = reset; // @[:@8874.4]
  assign S8DP1_6_io_int_in_A_0 = ff00_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@9053.4]
  assign S8DP1_6_io_int_in_A_1 = ff00_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@9054.4]
  assign S8DP1_6_io_int_in_A_2 = ff00_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@9055.4]
  assign S8DP1_6_io_int_in_A_3 = ff00_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@9056.4]
  assign S8DP1_6_io_int_in_A_4 = ff00_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@9057.4]
  assign S8DP1_6_io_int_in_A_5 = ff00_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@9058.4]
  assign S8DP1_6_io_int_in_A_6 = ff00_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@9059.4]
  assign S8DP1_6_io_int_in_A_7 = ff00_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@9060.4]
  assign S8DP1_6_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 55:21:@9052.4]
  assign S8DP1_6_io_tag_0 = ffb2_io_out_tag_2_0; // @[STA_VDBB.scala 55:21:@9044.4]
  assign S8DP1_6_io_tag_1 = ffb2_io_out_tag_2_1; // @[STA_VDBB.scala 55:21:@9045.4]
  assign S8DP1_6_io_tag_2 = ffb2_io_out_tag_2_2; // @[STA_VDBB.scala 55:21:@9046.4]
  assign S8DP1_6_io_tag_3 = ffb2_io_out_tag_2_3; // @[STA_VDBB.scala 55:21:@9047.4]
  assign S8DP1_6_io_tag_4 = ffb2_io_out_tag_2_4; // @[STA_VDBB.scala 55:21:@9048.4]
  assign S8DP1_6_io_tag_5 = ffb2_io_out_tag_2_5; // @[STA_VDBB.scala 55:21:@9049.4]
  assign S8DP1_6_io_tag_6 = ffb2_io_out_tag_2_6; // @[STA_VDBB.scala 55:21:@9050.4]
  assign S8DP1_6_io_tag_7 = ffb2_io_out_tag_2_7; // @[STA_VDBB.scala 55:21:@9051.4]
  assign S8DP1_7_clock = clock; // @[:@8876.4]
  assign S8DP1_7_reset = reset; // @[:@8877.4]
  assign S8DP1_7_io_int_in_A_0 = ff00_io_out_data_0_0; // @[STA_VDBB.scala 55:21:@9079.4]
  assign S8DP1_7_io_int_in_A_1 = ff00_io_out_data_0_1; // @[STA_VDBB.scala 55:21:@9080.4]
  assign S8DP1_7_io_int_in_A_2 = ff00_io_out_data_0_2; // @[STA_VDBB.scala 55:21:@9081.4]
  assign S8DP1_7_io_int_in_A_3 = ff00_io_out_data_0_3; // @[STA_VDBB.scala 55:21:@9082.4]
  assign S8DP1_7_io_int_in_A_4 = ff00_io_out_data_0_4; // @[STA_VDBB.scala 55:21:@9083.4]
  assign S8DP1_7_io_int_in_A_5 = ff00_io_out_data_0_5; // @[STA_VDBB.scala 55:21:@9084.4]
  assign S8DP1_7_io_int_in_A_6 = ff00_io_out_data_0_6; // @[STA_VDBB.scala 55:21:@9085.4]
  assign S8DP1_7_io_int_in_A_7 = ff00_io_out_data_0_7; // @[STA_VDBB.scala 55:21:@9086.4]
  assign S8DP1_7_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 55:21:@9078.4]
  assign S8DP1_7_io_tag_0 = ffb2_io_out_tag_3_0; // @[STA_VDBB.scala 55:21:@9070.4]
  assign S8DP1_7_io_tag_1 = ffb2_io_out_tag_3_1; // @[STA_VDBB.scala 55:21:@9071.4]
  assign S8DP1_7_io_tag_2 = ffb2_io_out_tag_3_2; // @[STA_VDBB.scala 55:21:@9072.4]
  assign S8DP1_7_io_tag_3 = ffb2_io_out_tag_3_3; // @[STA_VDBB.scala 55:21:@9073.4]
  assign S8DP1_7_io_tag_4 = ffb2_io_out_tag_3_4; // @[STA_VDBB.scala 55:21:@9074.4]
  assign S8DP1_7_io_tag_5 = ffb2_io_out_tag_3_5; // @[STA_VDBB.scala 55:21:@9075.4]
  assign S8DP1_7_io_tag_6 = ffb2_io_out_tag_3_6; // @[STA_VDBB.scala 55:21:@9076.4]
  assign S8DP1_7_io_tag_7 = ffb2_io_out_tag_3_7; // @[STA_VDBB.scala 55:21:@9077.4]
  assign S8DP1_8_clock = clock; // @[:@9088.4]
  assign S8DP1_8_reset = reset; // @[:@9089.4]
  assign S8DP1_8_io_int_in_A_0 = ffa1_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9130.4]
  assign S8DP1_8_io_int_in_A_1 = ffa1_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9131.4]
  assign S8DP1_8_io_int_in_A_2 = ffa1_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9132.4]
  assign S8DP1_8_io_int_in_A_3 = ffa1_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9133.4]
  assign S8DP1_8_io_int_in_A_4 = ffa1_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9134.4]
  assign S8DP1_8_io_int_in_A_5 = ffa1_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9135.4]
  assign S8DP1_8_io_int_in_A_6 = ffa1_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9136.4]
  assign S8DP1_8_io_int_in_A_7 = ffa1_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9137.4]
  assign S8DP1_8_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 56:21:@9129.4]
  assign S8DP1_8_io_tag_0 = ffb1_io_out_tag_0_0; // @[STA_VDBB.scala 56:21:@9121.4]
  assign S8DP1_8_io_tag_1 = ffb1_io_out_tag_0_1; // @[STA_VDBB.scala 56:21:@9122.4]
  assign S8DP1_8_io_tag_2 = ffb1_io_out_tag_0_2; // @[STA_VDBB.scala 56:21:@9123.4]
  assign S8DP1_8_io_tag_3 = ffb1_io_out_tag_0_3; // @[STA_VDBB.scala 56:21:@9124.4]
  assign S8DP1_8_io_tag_4 = ffb1_io_out_tag_0_4; // @[STA_VDBB.scala 56:21:@9125.4]
  assign S8DP1_8_io_tag_5 = ffb1_io_out_tag_0_5; // @[STA_VDBB.scala 56:21:@9126.4]
  assign S8DP1_8_io_tag_6 = ffb1_io_out_tag_0_6; // @[STA_VDBB.scala 56:21:@9127.4]
  assign S8DP1_8_io_tag_7 = ffb1_io_out_tag_0_7; // @[STA_VDBB.scala 56:21:@9128.4]
  assign S8DP1_9_clock = clock; // @[:@9091.4]
  assign S8DP1_9_reset = reset; // @[:@9092.4]
  assign S8DP1_9_io_int_in_A_0 = ffa1_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9156.4]
  assign S8DP1_9_io_int_in_A_1 = ffa1_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9157.4]
  assign S8DP1_9_io_int_in_A_2 = ffa1_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9158.4]
  assign S8DP1_9_io_int_in_A_3 = ffa1_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9159.4]
  assign S8DP1_9_io_int_in_A_4 = ffa1_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9160.4]
  assign S8DP1_9_io_int_in_A_5 = ffa1_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9161.4]
  assign S8DP1_9_io_int_in_A_6 = ffa1_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9162.4]
  assign S8DP1_9_io_int_in_A_7 = ffa1_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9163.4]
  assign S8DP1_9_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 56:21:@9155.4]
  assign S8DP1_9_io_tag_0 = ffb1_io_out_tag_1_0; // @[STA_VDBB.scala 56:21:@9147.4]
  assign S8DP1_9_io_tag_1 = ffb1_io_out_tag_1_1; // @[STA_VDBB.scala 56:21:@9148.4]
  assign S8DP1_9_io_tag_2 = ffb1_io_out_tag_1_2; // @[STA_VDBB.scala 56:21:@9149.4]
  assign S8DP1_9_io_tag_3 = ffb1_io_out_tag_1_3; // @[STA_VDBB.scala 56:21:@9150.4]
  assign S8DP1_9_io_tag_4 = ffb1_io_out_tag_1_4; // @[STA_VDBB.scala 56:21:@9151.4]
  assign S8DP1_9_io_tag_5 = ffb1_io_out_tag_1_5; // @[STA_VDBB.scala 56:21:@9152.4]
  assign S8DP1_9_io_tag_6 = ffb1_io_out_tag_1_6; // @[STA_VDBB.scala 56:21:@9153.4]
  assign S8DP1_9_io_tag_7 = ffb1_io_out_tag_1_7; // @[STA_VDBB.scala 56:21:@9154.4]
  assign S8DP1_10_clock = clock; // @[:@9094.4]
  assign S8DP1_10_reset = reset; // @[:@9095.4]
  assign S8DP1_10_io_int_in_A_0 = ffa1_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9182.4]
  assign S8DP1_10_io_int_in_A_1 = ffa1_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9183.4]
  assign S8DP1_10_io_int_in_A_2 = ffa1_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9184.4]
  assign S8DP1_10_io_int_in_A_3 = ffa1_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9185.4]
  assign S8DP1_10_io_int_in_A_4 = ffa1_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9186.4]
  assign S8DP1_10_io_int_in_A_5 = ffa1_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9187.4]
  assign S8DP1_10_io_int_in_A_6 = ffa1_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9188.4]
  assign S8DP1_10_io_int_in_A_7 = ffa1_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9189.4]
  assign S8DP1_10_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 56:21:@9181.4]
  assign S8DP1_10_io_tag_0 = ffb1_io_out_tag_2_0; // @[STA_VDBB.scala 56:21:@9173.4]
  assign S8DP1_10_io_tag_1 = ffb1_io_out_tag_2_1; // @[STA_VDBB.scala 56:21:@9174.4]
  assign S8DP1_10_io_tag_2 = ffb1_io_out_tag_2_2; // @[STA_VDBB.scala 56:21:@9175.4]
  assign S8DP1_10_io_tag_3 = ffb1_io_out_tag_2_3; // @[STA_VDBB.scala 56:21:@9176.4]
  assign S8DP1_10_io_tag_4 = ffb1_io_out_tag_2_4; // @[STA_VDBB.scala 56:21:@9177.4]
  assign S8DP1_10_io_tag_5 = ffb1_io_out_tag_2_5; // @[STA_VDBB.scala 56:21:@9178.4]
  assign S8DP1_10_io_tag_6 = ffb1_io_out_tag_2_6; // @[STA_VDBB.scala 56:21:@9179.4]
  assign S8DP1_10_io_tag_7 = ffb1_io_out_tag_2_7; // @[STA_VDBB.scala 56:21:@9180.4]
  assign S8DP1_11_clock = clock; // @[:@9097.4]
  assign S8DP1_11_reset = reset; // @[:@9098.4]
  assign S8DP1_11_io_int_in_A_0 = ffa1_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9208.4]
  assign S8DP1_11_io_int_in_A_1 = ffa1_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9209.4]
  assign S8DP1_11_io_int_in_A_2 = ffa1_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9210.4]
  assign S8DP1_11_io_int_in_A_3 = ffa1_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9211.4]
  assign S8DP1_11_io_int_in_A_4 = ffa1_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9212.4]
  assign S8DP1_11_io_int_in_A_5 = ffa1_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9213.4]
  assign S8DP1_11_io_int_in_A_6 = ffa1_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9214.4]
  assign S8DP1_11_io_int_in_A_7 = ffa1_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9215.4]
  assign S8DP1_11_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 56:21:@9207.4]
  assign S8DP1_11_io_tag_0 = ffb1_io_out_tag_3_0; // @[STA_VDBB.scala 56:21:@9199.4]
  assign S8DP1_11_io_tag_1 = ffb1_io_out_tag_3_1; // @[STA_VDBB.scala 56:21:@9200.4]
  assign S8DP1_11_io_tag_2 = ffb1_io_out_tag_3_2; // @[STA_VDBB.scala 56:21:@9201.4]
  assign S8DP1_11_io_tag_3 = ffb1_io_out_tag_3_3; // @[STA_VDBB.scala 56:21:@9202.4]
  assign S8DP1_11_io_tag_4 = ffb1_io_out_tag_3_4; // @[STA_VDBB.scala 56:21:@9203.4]
  assign S8DP1_11_io_tag_5 = ffb1_io_out_tag_3_5; // @[STA_VDBB.scala 56:21:@9204.4]
  assign S8DP1_11_io_tag_6 = ffb1_io_out_tag_3_6; // @[STA_VDBB.scala 56:21:@9205.4]
  assign S8DP1_11_io_tag_7 = ffb1_io_out_tag_3_7; // @[STA_VDBB.scala 56:21:@9206.4]
  assign S8DP1_12_clock = clock; // @[:@9100.4]
  assign S8DP1_12_reset = reset; // @[:@9101.4]
  assign S8DP1_12_io_int_in_A_0 = ff00_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9234.4]
  assign S8DP1_12_io_int_in_A_1 = ff00_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9235.4]
  assign S8DP1_12_io_int_in_A_2 = ff00_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9236.4]
  assign S8DP1_12_io_int_in_A_3 = ff00_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9237.4]
  assign S8DP1_12_io_int_in_A_4 = ff00_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9238.4]
  assign S8DP1_12_io_int_in_A_5 = ff00_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9239.4]
  assign S8DP1_12_io_int_in_A_6 = ff00_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9240.4]
  assign S8DP1_12_io_int_in_A_7 = ff00_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9241.4]
  assign S8DP1_12_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 56:21:@9233.4]
  assign S8DP1_12_io_tag_0 = ffb2_io_out_tag_0_0; // @[STA_VDBB.scala 56:21:@9225.4]
  assign S8DP1_12_io_tag_1 = ffb2_io_out_tag_0_1; // @[STA_VDBB.scala 56:21:@9226.4]
  assign S8DP1_12_io_tag_2 = ffb2_io_out_tag_0_2; // @[STA_VDBB.scala 56:21:@9227.4]
  assign S8DP1_12_io_tag_3 = ffb2_io_out_tag_0_3; // @[STA_VDBB.scala 56:21:@9228.4]
  assign S8DP1_12_io_tag_4 = ffb2_io_out_tag_0_4; // @[STA_VDBB.scala 56:21:@9229.4]
  assign S8DP1_12_io_tag_5 = ffb2_io_out_tag_0_5; // @[STA_VDBB.scala 56:21:@9230.4]
  assign S8DP1_12_io_tag_6 = ffb2_io_out_tag_0_6; // @[STA_VDBB.scala 56:21:@9231.4]
  assign S8DP1_12_io_tag_7 = ffb2_io_out_tag_0_7; // @[STA_VDBB.scala 56:21:@9232.4]
  assign S8DP1_13_clock = clock; // @[:@9103.4]
  assign S8DP1_13_reset = reset; // @[:@9104.4]
  assign S8DP1_13_io_int_in_A_0 = ff00_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9260.4]
  assign S8DP1_13_io_int_in_A_1 = ff00_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9261.4]
  assign S8DP1_13_io_int_in_A_2 = ff00_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9262.4]
  assign S8DP1_13_io_int_in_A_3 = ff00_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9263.4]
  assign S8DP1_13_io_int_in_A_4 = ff00_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9264.4]
  assign S8DP1_13_io_int_in_A_5 = ff00_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9265.4]
  assign S8DP1_13_io_int_in_A_6 = ff00_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9266.4]
  assign S8DP1_13_io_int_in_A_7 = ff00_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9267.4]
  assign S8DP1_13_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 56:21:@9259.4]
  assign S8DP1_13_io_tag_0 = ffb2_io_out_tag_1_0; // @[STA_VDBB.scala 56:21:@9251.4]
  assign S8DP1_13_io_tag_1 = ffb2_io_out_tag_1_1; // @[STA_VDBB.scala 56:21:@9252.4]
  assign S8DP1_13_io_tag_2 = ffb2_io_out_tag_1_2; // @[STA_VDBB.scala 56:21:@9253.4]
  assign S8DP1_13_io_tag_3 = ffb2_io_out_tag_1_3; // @[STA_VDBB.scala 56:21:@9254.4]
  assign S8DP1_13_io_tag_4 = ffb2_io_out_tag_1_4; // @[STA_VDBB.scala 56:21:@9255.4]
  assign S8DP1_13_io_tag_5 = ffb2_io_out_tag_1_5; // @[STA_VDBB.scala 56:21:@9256.4]
  assign S8DP1_13_io_tag_6 = ffb2_io_out_tag_1_6; // @[STA_VDBB.scala 56:21:@9257.4]
  assign S8DP1_13_io_tag_7 = ffb2_io_out_tag_1_7; // @[STA_VDBB.scala 56:21:@9258.4]
  assign S8DP1_14_clock = clock; // @[:@9106.4]
  assign S8DP1_14_reset = reset; // @[:@9107.4]
  assign S8DP1_14_io_int_in_A_0 = ff00_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9286.4]
  assign S8DP1_14_io_int_in_A_1 = ff00_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9287.4]
  assign S8DP1_14_io_int_in_A_2 = ff00_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9288.4]
  assign S8DP1_14_io_int_in_A_3 = ff00_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9289.4]
  assign S8DP1_14_io_int_in_A_4 = ff00_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9290.4]
  assign S8DP1_14_io_int_in_A_5 = ff00_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9291.4]
  assign S8DP1_14_io_int_in_A_6 = ff00_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9292.4]
  assign S8DP1_14_io_int_in_A_7 = ff00_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9293.4]
  assign S8DP1_14_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 56:21:@9285.4]
  assign S8DP1_14_io_tag_0 = ffb2_io_out_tag_2_0; // @[STA_VDBB.scala 56:21:@9277.4]
  assign S8DP1_14_io_tag_1 = ffb2_io_out_tag_2_1; // @[STA_VDBB.scala 56:21:@9278.4]
  assign S8DP1_14_io_tag_2 = ffb2_io_out_tag_2_2; // @[STA_VDBB.scala 56:21:@9279.4]
  assign S8DP1_14_io_tag_3 = ffb2_io_out_tag_2_3; // @[STA_VDBB.scala 56:21:@9280.4]
  assign S8DP1_14_io_tag_4 = ffb2_io_out_tag_2_4; // @[STA_VDBB.scala 56:21:@9281.4]
  assign S8DP1_14_io_tag_5 = ffb2_io_out_tag_2_5; // @[STA_VDBB.scala 56:21:@9282.4]
  assign S8DP1_14_io_tag_6 = ffb2_io_out_tag_2_6; // @[STA_VDBB.scala 56:21:@9283.4]
  assign S8DP1_14_io_tag_7 = ffb2_io_out_tag_2_7; // @[STA_VDBB.scala 56:21:@9284.4]
  assign S8DP1_15_clock = clock; // @[:@9109.4]
  assign S8DP1_15_reset = reset; // @[:@9110.4]
  assign S8DP1_15_io_int_in_A_0 = ff00_io_out_data_1_0; // @[STA_VDBB.scala 56:21:@9312.4]
  assign S8DP1_15_io_int_in_A_1 = ff00_io_out_data_1_1; // @[STA_VDBB.scala 56:21:@9313.4]
  assign S8DP1_15_io_int_in_A_2 = ff00_io_out_data_1_2; // @[STA_VDBB.scala 56:21:@9314.4]
  assign S8DP1_15_io_int_in_A_3 = ff00_io_out_data_1_3; // @[STA_VDBB.scala 56:21:@9315.4]
  assign S8DP1_15_io_int_in_A_4 = ff00_io_out_data_1_4; // @[STA_VDBB.scala 56:21:@9316.4]
  assign S8DP1_15_io_int_in_A_5 = ff00_io_out_data_1_5; // @[STA_VDBB.scala 56:21:@9317.4]
  assign S8DP1_15_io_int_in_A_6 = ff00_io_out_data_1_6; // @[STA_VDBB.scala 56:21:@9318.4]
  assign S8DP1_15_io_int_in_A_7 = ff00_io_out_data_1_7; // @[STA_VDBB.scala 56:21:@9319.4]
  assign S8DP1_15_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 56:21:@9311.4]
  assign S8DP1_15_io_tag_0 = ffb2_io_out_tag_3_0; // @[STA_VDBB.scala 56:21:@9303.4]
  assign S8DP1_15_io_tag_1 = ffb2_io_out_tag_3_1; // @[STA_VDBB.scala 56:21:@9304.4]
  assign S8DP1_15_io_tag_2 = ffb2_io_out_tag_3_2; // @[STA_VDBB.scala 56:21:@9305.4]
  assign S8DP1_15_io_tag_3 = ffb2_io_out_tag_3_3; // @[STA_VDBB.scala 56:21:@9306.4]
  assign S8DP1_15_io_tag_4 = ffb2_io_out_tag_3_4; // @[STA_VDBB.scala 56:21:@9307.4]
  assign S8DP1_15_io_tag_5 = ffb2_io_out_tag_3_5; // @[STA_VDBB.scala 56:21:@9308.4]
  assign S8DP1_15_io_tag_6 = ffb2_io_out_tag_3_6; // @[STA_VDBB.scala 56:21:@9309.4]
  assign S8DP1_15_io_tag_7 = ffb2_io_out_tag_3_7; // @[STA_VDBB.scala 56:21:@9310.4]
  assign S8DP1_16_clock = clock; // @[:@9321.4]
  assign S8DP1_16_reset = reset; // @[:@9322.4]
  assign S8DP1_16_io_int_in_A_0 = ff01_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9363.4]
  assign S8DP1_16_io_int_in_A_1 = ff01_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9364.4]
  assign S8DP1_16_io_int_in_A_2 = ff01_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9365.4]
  assign S8DP1_16_io_int_in_A_3 = ff01_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9366.4]
  assign S8DP1_16_io_int_in_A_4 = ff01_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9367.4]
  assign S8DP1_16_io_int_in_A_5 = ff01_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9368.4]
  assign S8DP1_16_io_int_in_A_6 = ff01_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9369.4]
  assign S8DP1_16_io_int_in_A_7 = ff01_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9370.4]
  assign S8DP1_16_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 57:21:@9362.4]
  assign S8DP1_16_io_tag_0 = ff01_io_out_tag_0_0; // @[STA_VDBB.scala 57:21:@9354.4]
  assign S8DP1_16_io_tag_1 = ff01_io_out_tag_0_1; // @[STA_VDBB.scala 57:21:@9355.4]
  assign S8DP1_16_io_tag_2 = ff01_io_out_tag_0_2; // @[STA_VDBB.scala 57:21:@9356.4]
  assign S8DP1_16_io_tag_3 = ff01_io_out_tag_0_3; // @[STA_VDBB.scala 57:21:@9357.4]
  assign S8DP1_16_io_tag_4 = ff01_io_out_tag_0_4; // @[STA_VDBB.scala 57:21:@9358.4]
  assign S8DP1_16_io_tag_5 = ff01_io_out_tag_0_5; // @[STA_VDBB.scala 57:21:@9359.4]
  assign S8DP1_16_io_tag_6 = ff01_io_out_tag_0_6; // @[STA_VDBB.scala 57:21:@9360.4]
  assign S8DP1_16_io_tag_7 = ff01_io_out_tag_0_7; // @[STA_VDBB.scala 57:21:@9361.4]
  assign S8DP1_17_clock = clock; // @[:@9324.4]
  assign S8DP1_17_reset = reset; // @[:@9325.4]
  assign S8DP1_17_io_int_in_A_0 = ff01_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9389.4]
  assign S8DP1_17_io_int_in_A_1 = ff01_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9390.4]
  assign S8DP1_17_io_int_in_A_2 = ff01_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9391.4]
  assign S8DP1_17_io_int_in_A_3 = ff01_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9392.4]
  assign S8DP1_17_io_int_in_A_4 = ff01_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9393.4]
  assign S8DP1_17_io_int_in_A_5 = ff01_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9394.4]
  assign S8DP1_17_io_int_in_A_6 = ff01_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9395.4]
  assign S8DP1_17_io_int_in_A_7 = ff01_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9396.4]
  assign S8DP1_17_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 57:21:@9388.4]
  assign S8DP1_17_io_tag_0 = ff01_io_out_tag_1_0; // @[STA_VDBB.scala 57:21:@9380.4]
  assign S8DP1_17_io_tag_1 = ff01_io_out_tag_1_1; // @[STA_VDBB.scala 57:21:@9381.4]
  assign S8DP1_17_io_tag_2 = ff01_io_out_tag_1_2; // @[STA_VDBB.scala 57:21:@9382.4]
  assign S8DP1_17_io_tag_3 = ff01_io_out_tag_1_3; // @[STA_VDBB.scala 57:21:@9383.4]
  assign S8DP1_17_io_tag_4 = ff01_io_out_tag_1_4; // @[STA_VDBB.scala 57:21:@9384.4]
  assign S8DP1_17_io_tag_5 = ff01_io_out_tag_1_5; // @[STA_VDBB.scala 57:21:@9385.4]
  assign S8DP1_17_io_tag_6 = ff01_io_out_tag_1_6; // @[STA_VDBB.scala 57:21:@9386.4]
  assign S8DP1_17_io_tag_7 = ff01_io_out_tag_1_7; // @[STA_VDBB.scala 57:21:@9387.4]
  assign S8DP1_18_clock = clock; // @[:@9327.4]
  assign S8DP1_18_reset = reset; // @[:@9328.4]
  assign S8DP1_18_io_int_in_A_0 = ff01_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9415.4]
  assign S8DP1_18_io_int_in_A_1 = ff01_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9416.4]
  assign S8DP1_18_io_int_in_A_2 = ff01_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9417.4]
  assign S8DP1_18_io_int_in_A_3 = ff01_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9418.4]
  assign S8DP1_18_io_int_in_A_4 = ff01_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9419.4]
  assign S8DP1_18_io_int_in_A_5 = ff01_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9420.4]
  assign S8DP1_18_io_int_in_A_6 = ff01_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9421.4]
  assign S8DP1_18_io_int_in_A_7 = ff01_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9422.4]
  assign S8DP1_18_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 57:21:@9414.4]
  assign S8DP1_18_io_tag_0 = ff01_io_out_tag_2_0; // @[STA_VDBB.scala 57:21:@9406.4]
  assign S8DP1_18_io_tag_1 = ff01_io_out_tag_2_1; // @[STA_VDBB.scala 57:21:@9407.4]
  assign S8DP1_18_io_tag_2 = ff01_io_out_tag_2_2; // @[STA_VDBB.scala 57:21:@9408.4]
  assign S8DP1_18_io_tag_3 = ff01_io_out_tag_2_3; // @[STA_VDBB.scala 57:21:@9409.4]
  assign S8DP1_18_io_tag_4 = ff01_io_out_tag_2_4; // @[STA_VDBB.scala 57:21:@9410.4]
  assign S8DP1_18_io_tag_5 = ff01_io_out_tag_2_5; // @[STA_VDBB.scala 57:21:@9411.4]
  assign S8DP1_18_io_tag_6 = ff01_io_out_tag_2_6; // @[STA_VDBB.scala 57:21:@9412.4]
  assign S8DP1_18_io_tag_7 = ff01_io_out_tag_2_7; // @[STA_VDBB.scala 57:21:@9413.4]
  assign S8DP1_19_clock = clock; // @[:@9330.4]
  assign S8DP1_19_reset = reset; // @[:@9331.4]
  assign S8DP1_19_io_int_in_A_0 = ff01_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9441.4]
  assign S8DP1_19_io_int_in_A_1 = ff01_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9442.4]
  assign S8DP1_19_io_int_in_A_2 = ff01_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9443.4]
  assign S8DP1_19_io_int_in_A_3 = ff01_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9444.4]
  assign S8DP1_19_io_int_in_A_4 = ff01_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9445.4]
  assign S8DP1_19_io_int_in_A_5 = ff01_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9446.4]
  assign S8DP1_19_io_int_in_A_6 = ff01_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9447.4]
  assign S8DP1_19_io_int_in_A_7 = ff01_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9448.4]
  assign S8DP1_19_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 57:21:@9440.4]
  assign S8DP1_19_io_tag_0 = ff01_io_out_tag_3_0; // @[STA_VDBB.scala 57:21:@9432.4]
  assign S8DP1_19_io_tag_1 = ff01_io_out_tag_3_1; // @[STA_VDBB.scala 57:21:@9433.4]
  assign S8DP1_19_io_tag_2 = ff01_io_out_tag_3_2; // @[STA_VDBB.scala 57:21:@9434.4]
  assign S8DP1_19_io_tag_3 = ff01_io_out_tag_3_3; // @[STA_VDBB.scala 57:21:@9435.4]
  assign S8DP1_19_io_tag_4 = ff01_io_out_tag_3_4; // @[STA_VDBB.scala 57:21:@9436.4]
  assign S8DP1_19_io_tag_5 = ff01_io_out_tag_3_5; // @[STA_VDBB.scala 57:21:@9437.4]
  assign S8DP1_19_io_tag_6 = ff01_io_out_tag_3_6; // @[STA_VDBB.scala 57:21:@9438.4]
  assign S8DP1_19_io_tag_7 = ff01_io_out_tag_3_7; // @[STA_VDBB.scala 57:21:@9439.4]
  assign S8DP1_20_clock = clock; // @[:@9333.4]
  assign S8DP1_20_reset = reset; // @[:@9334.4]
  assign S8DP1_20_io_int_in_A_0 = ff11_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9467.4]
  assign S8DP1_20_io_int_in_A_1 = ff11_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9468.4]
  assign S8DP1_20_io_int_in_A_2 = ff11_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9469.4]
  assign S8DP1_20_io_int_in_A_3 = ff11_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9470.4]
  assign S8DP1_20_io_int_in_A_4 = ff11_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9471.4]
  assign S8DP1_20_io_int_in_A_5 = ff11_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9472.4]
  assign S8DP1_20_io_int_in_A_6 = ff11_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9473.4]
  assign S8DP1_20_io_int_in_A_7 = ff11_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9474.4]
  assign S8DP1_20_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 57:21:@9466.4]
  assign S8DP1_20_io_tag_0 = ff10_io_out_tag_0_0; // @[STA_VDBB.scala 57:21:@9458.4]
  assign S8DP1_20_io_tag_1 = ff10_io_out_tag_0_1; // @[STA_VDBB.scala 57:21:@9459.4]
  assign S8DP1_20_io_tag_2 = ff10_io_out_tag_0_2; // @[STA_VDBB.scala 57:21:@9460.4]
  assign S8DP1_20_io_tag_3 = ff10_io_out_tag_0_3; // @[STA_VDBB.scala 57:21:@9461.4]
  assign S8DP1_20_io_tag_4 = ff10_io_out_tag_0_4; // @[STA_VDBB.scala 57:21:@9462.4]
  assign S8DP1_20_io_tag_5 = ff10_io_out_tag_0_5; // @[STA_VDBB.scala 57:21:@9463.4]
  assign S8DP1_20_io_tag_6 = ff10_io_out_tag_0_6; // @[STA_VDBB.scala 57:21:@9464.4]
  assign S8DP1_20_io_tag_7 = ff10_io_out_tag_0_7; // @[STA_VDBB.scala 57:21:@9465.4]
  assign S8DP1_21_clock = clock; // @[:@9336.4]
  assign S8DP1_21_reset = reset; // @[:@9337.4]
  assign S8DP1_21_io_int_in_A_0 = ff11_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9493.4]
  assign S8DP1_21_io_int_in_A_1 = ff11_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9494.4]
  assign S8DP1_21_io_int_in_A_2 = ff11_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9495.4]
  assign S8DP1_21_io_int_in_A_3 = ff11_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9496.4]
  assign S8DP1_21_io_int_in_A_4 = ff11_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9497.4]
  assign S8DP1_21_io_int_in_A_5 = ff11_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9498.4]
  assign S8DP1_21_io_int_in_A_6 = ff11_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9499.4]
  assign S8DP1_21_io_int_in_A_7 = ff11_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9500.4]
  assign S8DP1_21_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 57:21:@9492.4]
  assign S8DP1_21_io_tag_0 = ff10_io_out_tag_1_0; // @[STA_VDBB.scala 57:21:@9484.4]
  assign S8DP1_21_io_tag_1 = ff10_io_out_tag_1_1; // @[STA_VDBB.scala 57:21:@9485.4]
  assign S8DP1_21_io_tag_2 = ff10_io_out_tag_1_2; // @[STA_VDBB.scala 57:21:@9486.4]
  assign S8DP1_21_io_tag_3 = ff10_io_out_tag_1_3; // @[STA_VDBB.scala 57:21:@9487.4]
  assign S8DP1_21_io_tag_4 = ff10_io_out_tag_1_4; // @[STA_VDBB.scala 57:21:@9488.4]
  assign S8DP1_21_io_tag_5 = ff10_io_out_tag_1_5; // @[STA_VDBB.scala 57:21:@9489.4]
  assign S8DP1_21_io_tag_6 = ff10_io_out_tag_1_6; // @[STA_VDBB.scala 57:21:@9490.4]
  assign S8DP1_21_io_tag_7 = ff10_io_out_tag_1_7; // @[STA_VDBB.scala 57:21:@9491.4]
  assign S8DP1_22_clock = clock; // @[:@9339.4]
  assign S8DP1_22_reset = reset; // @[:@9340.4]
  assign S8DP1_22_io_int_in_A_0 = ff11_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9519.4]
  assign S8DP1_22_io_int_in_A_1 = ff11_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9520.4]
  assign S8DP1_22_io_int_in_A_2 = ff11_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9521.4]
  assign S8DP1_22_io_int_in_A_3 = ff11_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9522.4]
  assign S8DP1_22_io_int_in_A_4 = ff11_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9523.4]
  assign S8DP1_22_io_int_in_A_5 = ff11_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9524.4]
  assign S8DP1_22_io_int_in_A_6 = ff11_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9525.4]
  assign S8DP1_22_io_int_in_A_7 = ff11_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9526.4]
  assign S8DP1_22_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 57:21:@9518.4]
  assign S8DP1_22_io_tag_0 = ff10_io_out_tag_2_0; // @[STA_VDBB.scala 57:21:@9510.4]
  assign S8DP1_22_io_tag_1 = ff10_io_out_tag_2_1; // @[STA_VDBB.scala 57:21:@9511.4]
  assign S8DP1_22_io_tag_2 = ff10_io_out_tag_2_2; // @[STA_VDBB.scala 57:21:@9512.4]
  assign S8DP1_22_io_tag_3 = ff10_io_out_tag_2_3; // @[STA_VDBB.scala 57:21:@9513.4]
  assign S8DP1_22_io_tag_4 = ff10_io_out_tag_2_4; // @[STA_VDBB.scala 57:21:@9514.4]
  assign S8DP1_22_io_tag_5 = ff10_io_out_tag_2_5; // @[STA_VDBB.scala 57:21:@9515.4]
  assign S8DP1_22_io_tag_6 = ff10_io_out_tag_2_6; // @[STA_VDBB.scala 57:21:@9516.4]
  assign S8DP1_22_io_tag_7 = ff10_io_out_tag_2_7; // @[STA_VDBB.scala 57:21:@9517.4]
  assign S8DP1_23_clock = clock; // @[:@9342.4]
  assign S8DP1_23_reset = reset; // @[:@9343.4]
  assign S8DP1_23_io_int_in_A_0 = ff11_io_out_data_0_0; // @[STA_VDBB.scala 57:21:@9545.4]
  assign S8DP1_23_io_int_in_A_1 = ff11_io_out_data_0_1; // @[STA_VDBB.scala 57:21:@9546.4]
  assign S8DP1_23_io_int_in_A_2 = ff11_io_out_data_0_2; // @[STA_VDBB.scala 57:21:@9547.4]
  assign S8DP1_23_io_int_in_A_3 = ff11_io_out_data_0_3; // @[STA_VDBB.scala 57:21:@9548.4]
  assign S8DP1_23_io_int_in_A_4 = ff11_io_out_data_0_4; // @[STA_VDBB.scala 57:21:@9549.4]
  assign S8DP1_23_io_int_in_A_5 = ff11_io_out_data_0_5; // @[STA_VDBB.scala 57:21:@9550.4]
  assign S8DP1_23_io_int_in_A_6 = ff11_io_out_data_0_6; // @[STA_VDBB.scala 57:21:@9551.4]
  assign S8DP1_23_io_int_in_A_7 = ff11_io_out_data_0_7; // @[STA_VDBB.scala 57:21:@9552.4]
  assign S8DP1_23_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 57:21:@9544.4]
  assign S8DP1_23_io_tag_0 = ff10_io_out_tag_3_0; // @[STA_VDBB.scala 57:21:@9536.4]
  assign S8DP1_23_io_tag_1 = ff10_io_out_tag_3_1; // @[STA_VDBB.scala 57:21:@9537.4]
  assign S8DP1_23_io_tag_2 = ff10_io_out_tag_3_2; // @[STA_VDBB.scala 57:21:@9538.4]
  assign S8DP1_23_io_tag_3 = ff10_io_out_tag_3_3; // @[STA_VDBB.scala 57:21:@9539.4]
  assign S8DP1_23_io_tag_4 = ff10_io_out_tag_3_4; // @[STA_VDBB.scala 57:21:@9540.4]
  assign S8DP1_23_io_tag_5 = ff10_io_out_tag_3_5; // @[STA_VDBB.scala 57:21:@9541.4]
  assign S8DP1_23_io_tag_6 = ff10_io_out_tag_3_6; // @[STA_VDBB.scala 57:21:@9542.4]
  assign S8DP1_23_io_tag_7 = ff10_io_out_tag_3_7; // @[STA_VDBB.scala 57:21:@9543.4]
  assign S8DP1_24_clock = clock; // @[:@9554.4]
  assign S8DP1_24_reset = reset; // @[:@9555.4]
  assign S8DP1_24_io_int_in_A_0 = ff01_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9596.4]
  assign S8DP1_24_io_int_in_A_1 = ff01_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9597.4]
  assign S8DP1_24_io_int_in_A_2 = ff01_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9598.4]
  assign S8DP1_24_io_int_in_A_3 = ff01_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9599.4]
  assign S8DP1_24_io_int_in_A_4 = ff01_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9600.4]
  assign S8DP1_24_io_int_in_A_5 = ff01_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9601.4]
  assign S8DP1_24_io_int_in_A_6 = ff01_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9602.4]
  assign S8DP1_24_io_int_in_A_7 = ff01_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9603.4]
  assign S8DP1_24_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 58:21:@9595.4]
  assign S8DP1_24_io_tag_0 = ff01_io_out_tag_0_0; // @[STA_VDBB.scala 58:21:@9587.4]
  assign S8DP1_24_io_tag_1 = ff01_io_out_tag_0_1; // @[STA_VDBB.scala 58:21:@9588.4]
  assign S8DP1_24_io_tag_2 = ff01_io_out_tag_0_2; // @[STA_VDBB.scala 58:21:@9589.4]
  assign S8DP1_24_io_tag_3 = ff01_io_out_tag_0_3; // @[STA_VDBB.scala 58:21:@9590.4]
  assign S8DP1_24_io_tag_4 = ff01_io_out_tag_0_4; // @[STA_VDBB.scala 58:21:@9591.4]
  assign S8DP1_24_io_tag_5 = ff01_io_out_tag_0_5; // @[STA_VDBB.scala 58:21:@9592.4]
  assign S8DP1_24_io_tag_6 = ff01_io_out_tag_0_6; // @[STA_VDBB.scala 58:21:@9593.4]
  assign S8DP1_24_io_tag_7 = ff01_io_out_tag_0_7; // @[STA_VDBB.scala 58:21:@9594.4]
  assign S8DP1_25_clock = clock; // @[:@9557.4]
  assign S8DP1_25_reset = reset; // @[:@9558.4]
  assign S8DP1_25_io_int_in_A_0 = ff01_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9622.4]
  assign S8DP1_25_io_int_in_A_1 = ff01_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9623.4]
  assign S8DP1_25_io_int_in_A_2 = ff01_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9624.4]
  assign S8DP1_25_io_int_in_A_3 = ff01_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9625.4]
  assign S8DP1_25_io_int_in_A_4 = ff01_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9626.4]
  assign S8DP1_25_io_int_in_A_5 = ff01_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9627.4]
  assign S8DP1_25_io_int_in_A_6 = ff01_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9628.4]
  assign S8DP1_25_io_int_in_A_7 = ff01_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9629.4]
  assign S8DP1_25_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 58:21:@9621.4]
  assign S8DP1_25_io_tag_0 = ff01_io_out_tag_1_0; // @[STA_VDBB.scala 58:21:@9613.4]
  assign S8DP1_25_io_tag_1 = ff01_io_out_tag_1_1; // @[STA_VDBB.scala 58:21:@9614.4]
  assign S8DP1_25_io_tag_2 = ff01_io_out_tag_1_2; // @[STA_VDBB.scala 58:21:@9615.4]
  assign S8DP1_25_io_tag_3 = ff01_io_out_tag_1_3; // @[STA_VDBB.scala 58:21:@9616.4]
  assign S8DP1_25_io_tag_4 = ff01_io_out_tag_1_4; // @[STA_VDBB.scala 58:21:@9617.4]
  assign S8DP1_25_io_tag_5 = ff01_io_out_tag_1_5; // @[STA_VDBB.scala 58:21:@9618.4]
  assign S8DP1_25_io_tag_6 = ff01_io_out_tag_1_6; // @[STA_VDBB.scala 58:21:@9619.4]
  assign S8DP1_25_io_tag_7 = ff01_io_out_tag_1_7; // @[STA_VDBB.scala 58:21:@9620.4]
  assign S8DP1_26_clock = clock; // @[:@9560.4]
  assign S8DP1_26_reset = reset; // @[:@9561.4]
  assign S8DP1_26_io_int_in_A_0 = ff01_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9648.4]
  assign S8DP1_26_io_int_in_A_1 = ff01_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9649.4]
  assign S8DP1_26_io_int_in_A_2 = ff01_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9650.4]
  assign S8DP1_26_io_int_in_A_3 = ff01_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9651.4]
  assign S8DP1_26_io_int_in_A_4 = ff01_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9652.4]
  assign S8DP1_26_io_int_in_A_5 = ff01_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9653.4]
  assign S8DP1_26_io_int_in_A_6 = ff01_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9654.4]
  assign S8DP1_26_io_int_in_A_7 = ff01_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9655.4]
  assign S8DP1_26_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 58:21:@9647.4]
  assign S8DP1_26_io_tag_0 = ff01_io_out_tag_2_0; // @[STA_VDBB.scala 58:21:@9639.4]
  assign S8DP1_26_io_tag_1 = ff01_io_out_tag_2_1; // @[STA_VDBB.scala 58:21:@9640.4]
  assign S8DP1_26_io_tag_2 = ff01_io_out_tag_2_2; // @[STA_VDBB.scala 58:21:@9641.4]
  assign S8DP1_26_io_tag_3 = ff01_io_out_tag_2_3; // @[STA_VDBB.scala 58:21:@9642.4]
  assign S8DP1_26_io_tag_4 = ff01_io_out_tag_2_4; // @[STA_VDBB.scala 58:21:@9643.4]
  assign S8DP1_26_io_tag_5 = ff01_io_out_tag_2_5; // @[STA_VDBB.scala 58:21:@9644.4]
  assign S8DP1_26_io_tag_6 = ff01_io_out_tag_2_6; // @[STA_VDBB.scala 58:21:@9645.4]
  assign S8DP1_26_io_tag_7 = ff01_io_out_tag_2_7; // @[STA_VDBB.scala 58:21:@9646.4]
  assign S8DP1_27_clock = clock; // @[:@9563.4]
  assign S8DP1_27_reset = reset; // @[:@9564.4]
  assign S8DP1_27_io_int_in_A_0 = ff01_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9674.4]
  assign S8DP1_27_io_int_in_A_1 = ff01_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9675.4]
  assign S8DP1_27_io_int_in_A_2 = ff01_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9676.4]
  assign S8DP1_27_io_int_in_A_3 = ff01_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9677.4]
  assign S8DP1_27_io_int_in_A_4 = ff01_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9678.4]
  assign S8DP1_27_io_int_in_A_5 = ff01_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9679.4]
  assign S8DP1_27_io_int_in_A_6 = ff01_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9680.4]
  assign S8DP1_27_io_int_in_A_7 = ff01_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9681.4]
  assign S8DP1_27_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 58:21:@9673.4]
  assign S8DP1_27_io_tag_0 = ff01_io_out_tag_3_0; // @[STA_VDBB.scala 58:21:@9665.4]
  assign S8DP1_27_io_tag_1 = ff01_io_out_tag_3_1; // @[STA_VDBB.scala 58:21:@9666.4]
  assign S8DP1_27_io_tag_2 = ff01_io_out_tag_3_2; // @[STA_VDBB.scala 58:21:@9667.4]
  assign S8DP1_27_io_tag_3 = ff01_io_out_tag_3_3; // @[STA_VDBB.scala 58:21:@9668.4]
  assign S8DP1_27_io_tag_4 = ff01_io_out_tag_3_4; // @[STA_VDBB.scala 58:21:@9669.4]
  assign S8DP1_27_io_tag_5 = ff01_io_out_tag_3_5; // @[STA_VDBB.scala 58:21:@9670.4]
  assign S8DP1_27_io_tag_6 = ff01_io_out_tag_3_6; // @[STA_VDBB.scala 58:21:@9671.4]
  assign S8DP1_27_io_tag_7 = ff01_io_out_tag_3_7; // @[STA_VDBB.scala 58:21:@9672.4]
  assign S8DP1_28_clock = clock; // @[:@9566.4]
  assign S8DP1_28_reset = reset; // @[:@9567.4]
  assign S8DP1_28_io_int_in_A_0 = ff11_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9700.4]
  assign S8DP1_28_io_int_in_A_1 = ff11_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9701.4]
  assign S8DP1_28_io_int_in_A_2 = ff11_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9702.4]
  assign S8DP1_28_io_int_in_A_3 = ff11_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9703.4]
  assign S8DP1_28_io_int_in_A_4 = ff11_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9704.4]
  assign S8DP1_28_io_int_in_A_5 = ff11_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9705.4]
  assign S8DP1_28_io_int_in_A_6 = ff11_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9706.4]
  assign S8DP1_28_io_int_in_A_7 = ff11_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9707.4]
  assign S8DP1_28_io_int_in_B = MUX8_io_choice; // @[STA_VDBB.scala 58:21:@9699.4]
  assign S8DP1_28_io_tag_0 = ff10_io_out_tag_0_0; // @[STA_VDBB.scala 58:21:@9691.4]
  assign S8DP1_28_io_tag_1 = ff10_io_out_tag_0_1; // @[STA_VDBB.scala 58:21:@9692.4]
  assign S8DP1_28_io_tag_2 = ff10_io_out_tag_0_2; // @[STA_VDBB.scala 58:21:@9693.4]
  assign S8DP1_28_io_tag_3 = ff10_io_out_tag_0_3; // @[STA_VDBB.scala 58:21:@9694.4]
  assign S8DP1_28_io_tag_4 = ff10_io_out_tag_0_4; // @[STA_VDBB.scala 58:21:@9695.4]
  assign S8DP1_28_io_tag_5 = ff10_io_out_tag_0_5; // @[STA_VDBB.scala 58:21:@9696.4]
  assign S8DP1_28_io_tag_6 = ff10_io_out_tag_0_6; // @[STA_VDBB.scala 58:21:@9697.4]
  assign S8DP1_28_io_tag_7 = ff10_io_out_tag_0_7; // @[STA_VDBB.scala 58:21:@9698.4]
  assign S8DP1_29_clock = clock; // @[:@9569.4]
  assign S8DP1_29_reset = reset; // @[:@9570.4]
  assign S8DP1_29_io_int_in_A_0 = ff11_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9726.4]
  assign S8DP1_29_io_int_in_A_1 = ff11_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9727.4]
  assign S8DP1_29_io_int_in_A_2 = ff11_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9728.4]
  assign S8DP1_29_io_int_in_A_3 = ff11_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9729.4]
  assign S8DP1_29_io_int_in_A_4 = ff11_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9730.4]
  assign S8DP1_29_io_int_in_A_5 = ff11_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9731.4]
  assign S8DP1_29_io_int_in_A_6 = ff11_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9732.4]
  assign S8DP1_29_io_int_in_A_7 = ff11_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9733.4]
  assign S8DP1_29_io_int_in_B = MUX8_1_io_choice; // @[STA_VDBB.scala 58:21:@9725.4]
  assign S8DP1_29_io_tag_0 = ff10_io_out_tag_1_0; // @[STA_VDBB.scala 58:21:@9717.4]
  assign S8DP1_29_io_tag_1 = ff10_io_out_tag_1_1; // @[STA_VDBB.scala 58:21:@9718.4]
  assign S8DP1_29_io_tag_2 = ff10_io_out_tag_1_2; // @[STA_VDBB.scala 58:21:@9719.4]
  assign S8DP1_29_io_tag_3 = ff10_io_out_tag_1_3; // @[STA_VDBB.scala 58:21:@9720.4]
  assign S8DP1_29_io_tag_4 = ff10_io_out_tag_1_4; // @[STA_VDBB.scala 58:21:@9721.4]
  assign S8DP1_29_io_tag_5 = ff10_io_out_tag_1_5; // @[STA_VDBB.scala 58:21:@9722.4]
  assign S8DP1_29_io_tag_6 = ff10_io_out_tag_1_6; // @[STA_VDBB.scala 58:21:@9723.4]
  assign S8DP1_29_io_tag_7 = ff10_io_out_tag_1_7; // @[STA_VDBB.scala 58:21:@9724.4]
  assign S8DP1_30_clock = clock; // @[:@9572.4]
  assign S8DP1_30_reset = reset; // @[:@9573.4]
  assign S8DP1_30_io_int_in_A_0 = ff11_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9752.4]
  assign S8DP1_30_io_int_in_A_1 = ff11_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9753.4]
  assign S8DP1_30_io_int_in_A_2 = ff11_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9754.4]
  assign S8DP1_30_io_int_in_A_3 = ff11_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9755.4]
  assign S8DP1_30_io_int_in_A_4 = ff11_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9756.4]
  assign S8DP1_30_io_int_in_A_5 = ff11_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9757.4]
  assign S8DP1_30_io_int_in_A_6 = ff11_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9758.4]
  assign S8DP1_30_io_int_in_A_7 = ff11_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9759.4]
  assign S8DP1_30_io_int_in_B = MUX8_2_io_choice; // @[STA_VDBB.scala 58:21:@9751.4]
  assign S8DP1_30_io_tag_0 = ff10_io_out_tag_2_0; // @[STA_VDBB.scala 58:21:@9743.4]
  assign S8DP1_30_io_tag_1 = ff10_io_out_tag_2_1; // @[STA_VDBB.scala 58:21:@9744.4]
  assign S8DP1_30_io_tag_2 = ff10_io_out_tag_2_2; // @[STA_VDBB.scala 58:21:@9745.4]
  assign S8DP1_30_io_tag_3 = ff10_io_out_tag_2_3; // @[STA_VDBB.scala 58:21:@9746.4]
  assign S8DP1_30_io_tag_4 = ff10_io_out_tag_2_4; // @[STA_VDBB.scala 58:21:@9747.4]
  assign S8DP1_30_io_tag_5 = ff10_io_out_tag_2_5; // @[STA_VDBB.scala 58:21:@9748.4]
  assign S8DP1_30_io_tag_6 = ff10_io_out_tag_2_6; // @[STA_VDBB.scala 58:21:@9749.4]
  assign S8DP1_30_io_tag_7 = ff10_io_out_tag_2_7; // @[STA_VDBB.scala 58:21:@9750.4]
  assign S8DP1_31_clock = clock; // @[:@9575.4]
  assign S8DP1_31_reset = reset; // @[:@9576.4]
  assign S8DP1_31_io_int_in_A_0 = ff11_io_out_data_1_0; // @[STA_VDBB.scala 58:21:@9778.4]
  assign S8DP1_31_io_int_in_A_1 = ff11_io_out_data_1_1; // @[STA_VDBB.scala 58:21:@9779.4]
  assign S8DP1_31_io_int_in_A_2 = ff11_io_out_data_1_2; // @[STA_VDBB.scala 58:21:@9780.4]
  assign S8DP1_31_io_int_in_A_3 = ff11_io_out_data_1_3; // @[STA_VDBB.scala 58:21:@9781.4]
  assign S8DP1_31_io_int_in_A_4 = ff11_io_out_data_1_4; // @[STA_VDBB.scala 58:21:@9782.4]
  assign S8DP1_31_io_int_in_A_5 = ff11_io_out_data_1_5; // @[STA_VDBB.scala 58:21:@9783.4]
  assign S8DP1_31_io_int_in_A_6 = ff11_io_out_data_1_6; // @[STA_VDBB.scala 58:21:@9784.4]
  assign S8DP1_31_io_int_in_A_7 = ff11_io_out_data_1_7; // @[STA_VDBB.scala 58:21:@9785.4]
  assign S8DP1_31_io_int_in_B = MUX8_3_io_choice; // @[STA_VDBB.scala 58:21:@9777.4]
  assign S8DP1_31_io_tag_0 = ff10_io_out_tag_3_0; // @[STA_VDBB.scala 58:21:@9769.4]
  assign S8DP1_31_io_tag_1 = ff10_io_out_tag_3_1; // @[STA_VDBB.scala 58:21:@9770.4]
  assign S8DP1_31_io_tag_2 = ff10_io_out_tag_3_2; // @[STA_VDBB.scala 58:21:@9771.4]
  assign S8DP1_31_io_tag_3 = ff10_io_out_tag_3_3; // @[STA_VDBB.scala 58:21:@9772.4]
  assign S8DP1_31_io_tag_4 = ff10_io_out_tag_3_4; // @[STA_VDBB.scala 58:21:@9773.4]
  assign S8DP1_31_io_tag_5 = ff10_io_out_tag_3_5; // @[STA_VDBB.scala 58:21:@9774.4]
  assign S8DP1_31_io_tag_6 = ff10_io_out_tag_3_6; // @[STA_VDBB.scala 58:21:@9775.4]
  assign S8DP1_31_io_tag_7 = ff10_io_out_tag_3_7; // @[STA_VDBB.scala 58:21:@9776.4]
  assign ffb1_clock = clock; // @[:@9787.4]
  assign ffb1_reset = reset; // @[:@9788.4]
  assign ffb1_io_in_data_0_0 = io_in_B_0_8; // @[STA_VDBB.scala 99:29:@10080.4 STA_VDBB.scala 233:29:@18912.4]
  assign ffb1_io_in_data_0_1 = io_in_B_0_9; // @[STA_VDBB.scala 99:29:@10092.4 STA_VDBB.scala 233:29:@18924.4]
  assign ffb1_io_in_data_0_2 = io_in_B_0_10; // @[STA_VDBB.scala 99:29:@10104.4 STA_VDBB.scala 233:29:@18936.4]
  assign ffb1_io_in_data_0_3 = io_in_B_0_11; // @[STA_VDBB.scala 99:29:@10116.4 STA_VDBB.scala 233:29:@18948.4]
  assign ffb1_io_in_data_0_4 = io_in_B_0_12; // @[STA_VDBB.scala 99:29:@10128.4 STA_VDBB.scala 233:29:@18960.4]
  assign ffb1_io_in_data_0_5 = io_in_B_0_13; // @[STA_VDBB.scala 99:29:@10140.4 STA_VDBB.scala 233:29:@18972.4]
  assign ffb1_io_in_data_0_6 = io_in_B_0_14; // @[STA_VDBB.scala 99:29:@10152.4 STA_VDBB.scala 233:29:@18984.4]
  assign ffb1_io_in_data_0_7 = io_in_B_0_15; // @[STA_VDBB.scala 99:29:@10164.4 STA_VDBB.scala 233:29:@18996.4]
  assign ffb1_io_in_data_1_0 = io_in_B_1_8; // @[STA_VDBB.scala 99:29:@10082.4 STA_VDBB.scala 233:29:@18914.4]
  assign ffb1_io_in_data_1_1 = io_in_B_1_9; // @[STA_VDBB.scala 99:29:@10094.4 STA_VDBB.scala 233:29:@18926.4]
  assign ffb1_io_in_data_1_2 = io_in_B_1_10; // @[STA_VDBB.scala 99:29:@10106.4 STA_VDBB.scala 233:29:@18938.4]
  assign ffb1_io_in_data_1_3 = io_in_B_1_11; // @[STA_VDBB.scala 99:29:@10118.4 STA_VDBB.scala 233:29:@18950.4]
  assign ffb1_io_in_data_1_4 = io_in_B_1_12; // @[STA_VDBB.scala 99:29:@10130.4 STA_VDBB.scala 233:29:@18962.4]
  assign ffb1_io_in_data_1_5 = io_in_B_1_13; // @[STA_VDBB.scala 99:29:@10142.4 STA_VDBB.scala 233:29:@18974.4]
  assign ffb1_io_in_data_1_6 = io_in_B_1_14; // @[STA_VDBB.scala 99:29:@10154.4 STA_VDBB.scala 233:29:@18986.4]
  assign ffb1_io_in_data_1_7 = io_in_B_1_15; // @[STA_VDBB.scala 99:29:@10166.4 STA_VDBB.scala 233:29:@18998.4]
  assign ffb1_io_in_data_2_0 = io_in_B_2_8; // @[STA_VDBB.scala 99:29:@10084.4 STA_VDBB.scala 233:29:@18916.4]
  assign ffb1_io_in_data_2_1 = io_in_B_2_9; // @[STA_VDBB.scala 99:29:@10096.4 STA_VDBB.scala 233:29:@18928.4]
  assign ffb1_io_in_data_2_2 = io_in_B_2_10; // @[STA_VDBB.scala 99:29:@10108.4 STA_VDBB.scala 233:29:@18940.4]
  assign ffb1_io_in_data_2_3 = io_in_B_2_11; // @[STA_VDBB.scala 99:29:@10120.4 STA_VDBB.scala 233:29:@18952.4]
  assign ffb1_io_in_data_2_4 = io_in_B_2_12; // @[STA_VDBB.scala 99:29:@10132.4 STA_VDBB.scala 233:29:@18964.4]
  assign ffb1_io_in_data_2_5 = io_in_B_2_13; // @[STA_VDBB.scala 99:29:@10144.4 STA_VDBB.scala 233:29:@18976.4]
  assign ffb1_io_in_data_2_6 = io_in_B_2_14; // @[STA_VDBB.scala 99:29:@10156.4 STA_VDBB.scala 233:29:@18988.4]
  assign ffb1_io_in_data_2_7 = io_in_B_2_15; // @[STA_VDBB.scala 99:29:@10168.4 STA_VDBB.scala 233:29:@19000.4]
  assign ffb1_io_in_data_3_0 = io_in_B_3_8; // @[STA_VDBB.scala 99:29:@10086.4 STA_VDBB.scala 233:29:@18918.4]
  assign ffb1_io_in_data_3_1 = io_in_B_3_9; // @[STA_VDBB.scala 99:29:@10098.4 STA_VDBB.scala 233:29:@18930.4]
  assign ffb1_io_in_data_3_2 = io_in_B_3_10; // @[STA_VDBB.scala 99:29:@10110.4 STA_VDBB.scala 233:29:@18942.4]
  assign ffb1_io_in_data_3_3 = io_in_B_3_11; // @[STA_VDBB.scala 99:29:@10122.4 STA_VDBB.scala 233:29:@18954.4]
  assign ffb1_io_in_data_3_4 = io_in_B_3_12; // @[STA_VDBB.scala 99:29:@10134.4 STA_VDBB.scala 233:29:@18966.4]
  assign ffb1_io_in_data_3_5 = io_in_B_3_13; // @[STA_VDBB.scala 99:29:@10146.4 STA_VDBB.scala 233:29:@18978.4]
  assign ffb1_io_in_data_3_6 = io_in_B_3_14; // @[STA_VDBB.scala 99:29:@10158.4 STA_VDBB.scala 233:29:@18990.4]
  assign ffb1_io_in_data_3_7 = io_in_B_3_15; // @[STA_VDBB.scala 99:29:@10170.4 STA_VDBB.scala 233:29:@19002.4]
  assign ffb1_io_in_tag_0_0 = S8DP1_12_io_out_tag_0; // @[STA_VDBB.scala 108:23:@10180.4 STA_VDBB.scala 127:29:@10301.4 STA_VDBB.scala 127:29:@10326.4 STA_VDBB.scala 127:29:@10565.4 STA_VDBB.scala 127:29:@10590.4 STA_VDBB.scala 127:29:@10829.4 STA_VDBB.scala 127:29:@10854.4 STA_VDBB.scala 127:29:@11093.4 STA_VDBB.scala 127:29:@11118.4 STA_VDBB.scala 127:29:@11357.4 STA_VDBB.scala 127:29:@11382.4 STA_VDBB.scala 127:29:@11621.4 STA_VDBB.scala 127:29:@11646.4 STA_VDBB.scala 127:29:@11885.4 STA_VDBB.scala 127:29:@11910.4 STA_VDBB.scala 127:29:@12149.4 STA_VDBB.scala 127:29:@12174.4 STA_VDBB.scala 207:29:@13133.4 STA_VDBB.scala 207:29:@13158.4 STA_VDBB.scala 207:29:@13925.4 STA_VDBB.scala 207:29:@13950.4 STA_VDBB.scala 207:29:@14717.4 STA_VDBB.scala 207:29:@14742.4 STA_VDBB.scala 207:29:@15509.4 STA_VDBB.scala 207:29:@15534.4 STA_VDBB.scala 207:29:@16301.4 STA_VDBB.scala 207:29:@16326.4 STA_VDBB.scala 207:29:@17093.4 STA_VDBB.scala 207:29:@17118.4 STA_VDBB.scala 207:29:@17885.4 STA_VDBB.scala 207:29:@17910.4 STA_VDBB.scala 207:29:@18677.4 STA_VDBB.scala 207:29:@18702.4 STA_VDBB.scala 241:23:@19012.4 STA_VDBB.scala 260:29:@19133.4 STA_VDBB.scala 260:29:@19158.4 STA_VDBB.scala 260:29:@19397.4 STA_VDBB.scala 260:29:@19422.4 STA_VDBB.scala 260:29:@19661.4 STA_VDBB.scala 260:29:@19686.4 STA_VDBB.scala 260:29:@19925.4 STA_VDBB.scala 260:29:@19950.4 STA_VDBB.scala 260:29:@20189.4 STA_VDBB.scala 260:29:@20214.4 STA_VDBB.scala 260:29:@20453.4 STA_VDBB.scala 260:29:@20478.4 STA_VDBB.scala 260:29:@20717.4 STA_VDBB.scala 260:29:@20742.4 STA_VDBB.scala 260:29:@20981.4 STA_VDBB.scala 260:29:@21006.4 STA_VDBB.scala 339:29:@21965.4 STA_VDBB.scala 339:29:@21990.4 STA_VDBB.scala 339:29:@22757.4 STA_VDBB.scala 339:29:@22782.4 STA_VDBB.scala 339:29:@23549.4 STA_VDBB.scala 339:29:@23574.4 STA_VDBB.scala 339:29:@24341.4 STA_VDBB.scala 339:29:@24366.4 STA_VDBB.scala 339:29:@25133.4 STA_VDBB.scala 339:29:@25158.4 STA_VDBB.scala 339:29:@25925.4 STA_VDBB.scala 339:29:@25950.4 STA_VDBB.scala 339:29:@26717.4 STA_VDBB.scala 339:29:@26742.4 STA_VDBB.scala 339:29:@27509.4 STA_VDBB.scala 339:29:@27534.4]
  assign ffb1_io_in_tag_0_1 = S8DP1_12_io_out_tag_1; // @[STA_VDBB.scala 108:23:@10181.4 STA_VDBB.scala 127:29:@10302.4 STA_VDBB.scala 127:29:@10327.4 STA_VDBB.scala 127:29:@10566.4 STA_VDBB.scala 127:29:@10591.4 STA_VDBB.scala 127:29:@10830.4 STA_VDBB.scala 127:29:@10855.4 STA_VDBB.scala 127:29:@11094.4 STA_VDBB.scala 127:29:@11119.4 STA_VDBB.scala 127:29:@11358.4 STA_VDBB.scala 127:29:@11383.4 STA_VDBB.scala 127:29:@11622.4 STA_VDBB.scala 127:29:@11647.4 STA_VDBB.scala 127:29:@11886.4 STA_VDBB.scala 127:29:@11911.4 STA_VDBB.scala 127:29:@12150.4 STA_VDBB.scala 127:29:@12175.4 STA_VDBB.scala 207:29:@13134.4 STA_VDBB.scala 207:29:@13159.4 STA_VDBB.scala 207:29:@13926.4 STA_VDBB.scala 207:29:@13951.4 STA_VDBB.scala 207:29:@14718.4 STA_VDBB.scala 207:29:@14743.4 STA_VDBB.scala 207:29:@15510.4 STA_VDBB.scala 207:29:@15535.4 STA_VDBB.scala 207:29:@16302.4 STA_VDBB.scala 207:29:@16327.4 STA_VDBB.scala 207:29:@17094.4 STA_VDBB.scala 207:29:@17119.4 STA_VDBB.scala 207:29:@17886.4 STA_VDBB.scala 207:29:@17911.4 STA_VDBB.scala 207:29:@18678.4 STA_VDBB.scala 207:29:@18703.4 STA_VDBB.scala 241:23:@19013.4 STA_VDBB.scala 260:29:@19134.4 STA_VDBB.scala 260:29:@19159.4 STA_VDBB.scala 260:29:@19398.4 STA_VDBB.scala 260:29:@19423.4 STA_VDBB.scala 260:29:@19662.4 STA_VDBB.scala 260:29:@19687.4 STA_VDBB.scala 260:29:@19926.4 STA_VDBB.scala 260:29:@19951.4 STA_VDBB.scala 260:29:@20190.4 STA_VDBB.scala 260:29:@20215.4 STA_VDBB.scala 260:29:@20454.4 STA_VDBB.scala 260:29:@20479.4 STA_VDBB.scala 260:29:@20718.4 STA_VDBB.scala 260:29:@20743.4 STA_VDBB.scala 260:29:@20982.4 STA_VDBB.scala 260:29:@21007.4 STA_VDBB.scala 339:29:@21966.4 STA_VDBB.scala 339:29:@21991.4 STA_VDBB.scala 339:29:@22758.4 STA_VDBB.scala 339:29:@22783.4 STA_VDBB.scala 339:29:@23550.4 STA_VDBB.scala 339:29:@23575.4 STA_VDBB.scala 339:29:@24342.4 STA_VDBB.scala 339:29:@24367.4 STA_VDBB.scala 339:29:@25134.4 STA_VDBB.scala 339:29:@25159.4 STA_VDBB.scala 339:29:@25926.4 STA_VDBB.scala 339:29:@25951.4 STA_VDBB.scala 339:29:@26718.4 STA_VDBB.scala 339:29:@26743.4 STA_VDBB.scala 339:29:@27510.4 STA_VDBB.scala 339:29:@27535.4]
  assign ffb1_io_in_tag_0_2 = S8DP1_12_io_out_tag_2; // @[STA_VDBB.scala 108:23:@10182.4 STA_VDBB.scala 127:29:@10303.4 STA_VDBB.scala 127:29:@10328.4 STA_VDBB.scala 127:29:@10567.4 STA_VDBB.scala 127:29:@10592.4 STA_VDBB.scala 127:29:@10831.4 STA_VDBB.scala 127:29:@10856.4 STA_VDBB.scala 127:29:@11095.4 STA_VDBB.scala 127:29:@11120.4 STA_VDBB.scala 127:29:@11359.4 STA_VDBB.scala 127:29:@11384.4 STA_VDBB.scala 127:29:@11623.4 STA_VDBB.scala 127:29:@11648.4 STA_VDBB.scala 127:29:@11887.4 STA_VDBB.scala 127:29:@11912.4 STA_VDBB.scala 127:29:@12151.4 STA_VDBB.scala 127:29:@12176.4 STA_VDBB.scala 207:29:@13135.4 STA_VDBB.scala 207:29:@13160.4 STA_VDBB.scala 207:29:@13927.4 STA_VDBB.scala 207:29:@13952.4 STA_VDBB.scala 207:29:@14719.4 STA_VDBB.scala 207:29:@14744.4 STA_VDBB.scala 207:29:@15511.4 STA_VDBB.scala 207:29:@15536.4 STA_VDBB.scala 207:29:@16303.4 STA_VDBB.scala 207:29:@16328.4 STA_VDBB.scala 207:29:@17095.4 STA_VDBB.scala 207:29:@17120.4 STA_VDBB.scala 207:29:@17887.4 STA_VDBB.scala 207:29:@17912.4 STA_VDBB.scala 207:29:@18679.4 STA_VDBB.scala 207:29:@18704.4 STA_VDBB.scala 241:23:@19014.4 STA_VDBB.scala 260:29:@19135.4 STA_VDBB.scala 260:29:@19160.4 STA_VDBB.scala 260:29:@19399.4 STA_VDBB.scala 260:29:@19424.4 STA_VDBB.scala 260:29:@19663.4 STA_VDBB.scala 260:29:@19688.4 STA_VDBB.scala 260:29:@19927.4 STA_VDBB.scala 260:29:@19952.4 STA_VDBB.scala 260:29:@20191.4 STA_VDBB.scala 260:29:@20216.4 STA_VDBB.scala 260:29:@20455.4 STA_VDBB.scala 260:29:@20480.4 STA_VDBB.scala 260:29:@20719.4 STA_VDBB.scala 260:29:@20744.4 STA_VDBB.scala 260:29:@20983.4 STA_VDBB.scala 260:29:@21008.4 STA_VDBB.scala 339:29:@21967.4 STA_VDBB.scala 339:29:@21992.4 STA_VDBB.scala 339:29:@22759.4 STA_VDBB.scala 339:29:@22784.4 STA_VDBB.scala 339:29:@23551.4 STA_VDBB.scala 339:29:@23576.4 STA_VDBB.scala 339:29:@24343.4 STA_VDBB.scala 339:29:@24368.4 STA_VDBB.scala 339:29:@25135.4 STA_VDBB.scala 339:29:@25160.4 STA_VDBB.scala 339:29:@25927.4 STA_VDBB.scala 339:29:@25952.4 STA_VDBB.scala 339:29:@26719.4 STA_VDBB.scala 339:29:@26744.4 STA_VDBB.scala 339:29:@27511.4 STA_VDBB.scala 339:29:@27536.4]
  assign ffb1_io_in_tag_0_3 = S8DP1_12_io_out_tag_3; // @[STA_VDBB.scala 108:23:@10183.4 STA_VDBB.scala 127:29:@10304.4 STA_VDBB.scala 127:29:@10329.4 STA_VDBB.scala 127:29:@10568.4 STA_VDBB.scala 127:29:@10593.4 STA_VDBB.scala 127:29:@10832.4 STA_VDBB.scala 127:29:@10857.4 STA_VDBB.scala 127:29:@11096.4 STA_VDBB.scala 127:29:@11121.4 STA_VDBB.scala 127:29:@11360.4 STA_VDBB.scala 127:29:@11385.4 STA_VDBB.scala 127:29:@11624.4 STA_VDBB.scala 127:29:@11649.4 STA_VDBB.scala 127:29:@11888.4 STA_VDBB.scala 127:29:@11913.4 STA_VDBB.scala 127:29:@12152.4 STA_VDBB.scala 127:29:@12177.4 STA_VDBB.scala 207:29:@13136.4 STA_VDBB.scala 207:29:@13161.4 STA_VDBB.scala 207:29:@13928.4 STA_VDBB.scala 207:29:@13953.4 STA_VDBB.scala 207:29:@14720.4 STA_VDBB.scala 207:29:@14745.4 STA_VDBB.scala 207:29:@15512.4 STA_VDBB.scala 207:29:@15537.4 STA_VDBB.scala 207:29:@16304.4 STA_VDBB.scala 207:29:@16329.4 STA_VDBB.scala 207:29:@17096.4 STA_VDBB.scala 207:29:@17121.4 STA_VDBB.scala 207:29:@17888.4 STA_VDBB.scala 207:29:@17913.4 STA_VDBB.scala 207:29:@18680.4 STA_VDBB.scala 207:29:@18705.4 STA_VDBB.scala 241:23:@19015.4 STA_VDBB.scala 260:29:@19136.4 STA_VDBB.scala 260:29:@19161.4 STA_VDBB.scala 260:29:@19400.4 STA_VDBB.scala 260:29:@19425.4 STA_VDBB.scala 260:29:@19664.4 STA_VDBB.scala 260:29:@19689.4 STA_VDBB.scala 260:29:@19928.4 STA_VDBB.scala 260:29:@19953.4 STA_VDBB.scala 260:29:@20192.4 STA_VDBB.scala 260:29:@20217.4 STA_VDBB.scala 260:29:@20456.4 STA_VDBB.scala 260:29:@20481.4 STA_VDBB.scala 260:29:@20720.4 STA_VDBB.scala 260:29:@20745.4 STA_VDBB.scala 260:29:@20984.4 STA_VDBB.scala 260:29:@21009.4 STA_VDBB.scala 339:29:@21968.4 STA_VDBB.scala 339:29:@21993.4 STA_VDBB.scala 339:29:@22760.4 STA_VDBB.scala 339:29:@22785.4 STA_VDBB.scala 339:29:@23552.4 STA_VDBB.scala 339:29:@23577.4 STA_VDBB.scala 339:29:@24344.4 STA_VDBB.scala 339:29:@24369.4 STA_VDBB.scala 339:29:@25136.4 STA_VDBB.scala 339:29:@25161.4 STA_VDBB.scala 339:29:@25928.4 STA_VDBB.scala 339:29:@25953.4 STA_VDBB.scala 339:29:@26720.4 STA_VDBB.scala 339:29:@26745.4 STA_VDBB.scala 339:29:@27512.4 STA_VDBB.scala 339:29:@27537.4]
  assign ffb1_io_in_tag_0_4 = S8DP1_12_io_out_tag_4; // @[STA_VDBB.scala 108:23:@10184.4 STA_VDBB.scala 127:29:@10305.4 STA_VDBB.scala 127:29:@10330.4 STA_VDBB.scala 127:29:@10569.4 STA_VDBB.scala 127:29:@10594.4 STA_VDBB.scala 127:29:@10833.4 STA_VDBB.scala 127:29:@10858.4 STA_VDBB.scala 127:29:@11097.4 STA_VDBB.scala 127:29:@11122.4 STA_VDBB.scala 127:29:@11361.4 STA_VDBB.scala 127:29:@11386.4 STA_VDBB.scala 127:29:@11625.4 STA_VDBB.scala 127:29:@11650.4 STA_VDBB.scala 127:29:@11889.4 STA_VDBB.scala 127:29:@11914.4 STA_VDBB.scala 127:29:@12153.4 STA_VDBB.scala 127:29:@12178.4 STA_VDBB.scala 207:29:@13137.4 STA_VDBB.scala 207:29:@13162.4 STA_VDBB.scala 207:29:@13929.4 STA_VDBB.scala 207:29:@13954.4 STA_VDBB.scala 207:29:@14721.4 STA_VDBB.scala 207:29:@14746.4 STA_VDBB.scala 207:29:@15513.4 STA_VDBB.scala 207:29:@15538.4 STA_VDBB.scala 207:29:@16305.4 STA_VDBB.scala 207:29:@16330.4 STA_VDBB.scala 207:29:@17097.4 STA_VDBB.scala 207:29:@17122.4 STA_VDBB.scala 207:29:@17889.4 STA_VDBB.scala 207:29:@17914.4 STA_VDBB.scala 207:29:@18681.4 STA_VDBB.scala 207:29:@18706.4 STA_VDBB.scala 241:23:@19016.4 STA_VDBB.scala 260:29:@19137.4 STA_VDBB.scala 260:29:@19162.4 STA_VDBB.scala 260:29:@19401.4 STA_VDBB.scala 260:29:@19426.4 STA_VDBB.scala 260:29:@19665.4 STA_VDBB.scala 260:29:@19690.4 STA_VDBB.scala 260:29:@19929.4 STA_VDBB.scala 260:29:@19954.4 STA_VDBB.scala 260:29:@20193.4 STA_VDBB.scala 260:29:@20218.4 STA_VDBB.scala 260:29:@20457.4 STA_VDBB.scala 260:29:@20482.4 STA_VDBB.scala 260:29:@20721.4 STA_VDBB.scala 260:29:@20746.4 STA_VDBB.scala 260:29:@20985.4 STA_VDBB.scala 260:29:@21010.4 STA_VDBB.scala 339:29:@21969.4 STA_VDBB.scala 339:29:@21994.4 STA_VDBB.scala 339:29:@22761.4 STA_VDBB.scala 339:29:@22786.4 STA_VDBB.scala 339:29:@23553.4 STA_VDBB.scala 339:29:@23578.4 STA_VDBB.scala 339:29:@24345.4 STA_VDBB.scala 339:29:@24370.4 STA_VDBB.scala 339:29:@25137.4 STA_VDBB.scala 339:29:@25162.4 STA_VDBB.scala 339:29:@25929.4 STA_VDBB.scala 339:29:@25954.4 STA_VDBB.scala 339:29:@26721.4 STA_VDBB.scala 339:29:@26746.4 STA_VDBB.scala 339:29:@27513.4 STA_VDBB.scala 339:29:@27538.4]
  assign ffb1_io_in_tag_0_5 = S8DP1_12_io_out_tag_5; // @[STA_VDBB.scala 108:23:@10185.4 STA_VDBB.scala 127:29:@10306.4 STA_VDBB.scala 127:29:@10331.4 STA_VDBB.scala 127:29:@10570.4 STA_VDBB.scala 127:29:@10595.4 STA_VDBB.scala 127:29:@10834.4 STA_VDBB.scala 127:29:@10859.4 STA_VDBB.scala 127:29:@11098.4 STA_VDBB.scala 127:29:@11123.4 STA_VDBB.scala 127:29:@11362.4 STA_VDBB.scala 127:29:@11387.4 STA_VDBB.scala 127:29:@11626.4 STA_VDBB.scala 127:29:@11651.4 STA_VDBB.scala 127:29:@11890.4 STA_VDBB.scala 127:29:@11915.4 STA_VDBB.scala 127:29:@12154.4 STA_VDBB.scala 127:29:@12179.4 STA_VDBB.scala 207:29:@13138.4 STA_VDBB.scala 207:29:@13163.4 STA_VDBB.scala 207:29:@13930.4 STA_VDBB.scala 207:29:@13955.4 STA_VDBB.scala 207:29:@14722.4 STA_VDBB.scala 207:29:@14747.4 STA_VDBB.scala 207:29:@15514.4 STA_VDBB.scala 207:29:@15539.4 STA_VDBB.scala 207:29:@16306.4 STA_VDBB.scala 207:29:@16331.4 STA_VDBB.scala 207:29:@17098.4 STA_VDBB.scala 207:29:@17123.4 STA_VDBB.scala 207:29:@17890.4 STA_VDBB.scala 207:29:@17915.4 STA_VDBB.scala 207:29:@18682.4 STA_VDBB.scala 207:29:@18707.4 STA_VDBB.scala 241:23:@19017.4 STA_VDBB.scala 260:29:@19138.4 STA_VDBB.scala 260:29:@19163.4 STA_VDBB.scala 260:29:@19402.4 STA_VDBB.scala 260:29:@19427.4 STA_VDBB.scala 260:29:@19666.4 STA_VDBB.scala 260:29:@19691.4 STA_VDBB.scala 260:29:@19930.4 STA_VDBB.scala 260:29:@19955.4 STA_VDBB.scala 260:29:@20194.4 STA_VDBB.scala 260:29:@20219.4 STA_VDBB.scala 260:29:@20458.4 STA_VDBB.scala 260:29:@20483.4 STA_VDBB.scala 260:29:@20722.4 STA_VDBB.scala 260:29:@20747.4 STA_VDBB.scala 260:29:@20986.4 STA_VDBB.scala 260:29:@21011.4 STA_VDBB.scala 339:29:@21970.4 STA_VDBB.scala 339:29:@21995.4 STA_VDBB.scala 339:29:@22762.4 STA_VDBB.scala 339:29:@22787.4 STA_VDBB.scala 339:29:@23554.4 STA_VDBB.scala 339:29:@23579.4 STA_VDBB.scala 339:29:@24346.4 STA_VDBB.scala 339:29:@24371.4 STA_VDBB.scala 339:29:@25138.4 STA_VDBB.scala 339:29:@25163.4 STA_VDBB.scala 339:29:@25930.4 STA_VDBB.scala 339:29:@25955.4 STA_VDBB.scala 339:29:@26722.4 STA_VDBB.scala 339:29:@26747.4 STA_VDBB.scala 339:29:@27514.4 STA_VDBB.scala 339:29:@27539.4]
  assign ffb1_io_in_tag_0_6 = S8DP1_12_io_out_tag_6; // @[STA_VDBB.scala 108:23:@10186.4 STA_VDBB.scala 127:29:@10307.4 STA_VDBB.scala 127:29:@10332.4 STA_VDBB.scala 127:29:@10571.4 STA_VDBB.scala 127:29:@10596.4 STA_VDBB.scala 127:29:@10835.4 STA_VDBB.scala 127:29:@10860.4 STA_VDBB.scala 127:29:@11099.4 STA_VDBB.scala 127:29:@11124.4 STA_VDBB.scala 127:29:@11363.4 STA_VDBB.scala 127:29:@11388.4 STA_VDBB.scala 127:29:@11627.4 STA_VDBB.scala 127:29:@11652.4 STA_VDBB.scala 127:29:@11891.4 STA_VDBB.scala 127:29:@11916.4 STA_VDBB.scala 127:29:@12155.4 STA_VDBB.scala 127:29:@12180.4 STA_VDBB.scala 207:29:@13139.4 STA_VDBB.scala 207:29:@13164.4 STA_VDBB.scala 207:29:@13931.4 STA_VDBB.scala 207:29:@13956.4 STA_VDBB.scala 207:29:@14723.4 STA_VDBB.scala 207:29:@14748.4 STA_VDBB.scala 207:29:@15515.4 STA_VDBB.scala 207:29:@15540.4 STA_VDBB.scala 207:29:@16307.4 STA_VDBB.scala 207:29:@16332.4 STA_VDBB.scala 207:29:@17099.4 STA_VDBB.scala 207:29:@17124.4 STA_VDBB.scala 207:29:@17891.4 STA_VDBB.scala 207:29:@17916.4 STA_VDBB.scala 207:29:@18683.4 STA_VDBB.scala 207:29:@18708.4 STA_VDBB.scala 241:23:@19018.4 STA_VDBB.scala 260:29:@19139.4 STA_VDBB.scala 260:29:@19164.4 STA_VDBB.scala 260:29:@19403.4 STA_VDBB.scala 260:29:@19428.4 STA_VDBB.scala 260:29:@19667.4 STA_VDBB.scala 260:29:@19692.4 STA_VDBB.scala 260:29:@19931.4 STA_VDBB.scala 260:29:@19956.4 STA_VDBB.scala 260:29:@20195.4 STA_VDBB.scala 260:29:@20220.4 STA_VDBB.scala 260:29:@20459.4 STA_VDBB.scala 260:29:@20484.4 STA_VDBB.scala 260:29:@20723.4 STA_VDBB.scala 260:29:@20748.4 STA_VDBB.scala 260:29:@20987.4 STA_VDBB.scala 260:29:@21012.4 STA_VDBB.scala 339:29:@21971.4 STA_VDBB.scala 339:29:@21996.4 STA_VDBB.scala 339:29:@22763.4 STA_VDBB.scala 339:29:@22788.4 STA_VDBB.scala 339:29:@23555.4 STA_VDBB.scala 339:29:@23580.4 STA_VDBB.scala 339:29:@24347.4 STA_VDBB.scala 339:29:@24372.4 STA_VDBB.scala 339:29:@25139.4 STA_VDBB.scala 339:29:@25164.4 STA_VDBB.scala 339:29:@25931.4 STA_VDBB.scala 339:29:@25956.4 STA_VDBB.scala 339:29:@26723.4 STA_VDBB.scala 339:29:@26748.4 STA_VDBB.scala 339:29:@27515.4 STA_VDBB.scala 339:29:@27540.4]
  assign ffb1_io_in_tag_0_7 = S8DP1_12_io_out_tag_7; // @[STA_VDBB.scala 108:23:@10187.4 STA_VDBB.scala 127:29:@10308.4 STA_VDBB.scala 127:29:@10333.4 STA_VDBB.scala 127:29:@10572.4 STA_VDBB.scala 127:29:@10597.4 STA_VDBB.scala 127:29:@10836.4 STA_VDBB.scala 127:29:@10861.4 STA_VDBB.scala 127:29:@11100.4 STA_VDBB.scala 127:29:@11125.4 STA_VDBB.scala 127:29:@11364.4 STA_VDBB.scala 127:29:@11389.4 STA_VDBB.scala 127:29:@11628.4 STA_VDBB.scala 127:29:@11653.4 STA_VDBB.scala 127:29:@11892.4 STA_VDBB.scala 127:29:@11917.4 STA_VDBB.scala 127:29:@12156.4 STA_VDBB.scala 127:29:@12181.4 STA_VDBB.scala 207:29:@13140.4 STA_VDBB.scala 207:29:@13165.4 STA_VDBB.scala 207:29:@13932.4 STA_VDBB.scala 207:29:@13957.4 STA_VDBB.scala 207:29:@14724.4 STA_VDBB.scala 207:29:@14749.4 STA_VDBB.scala 207:29:@15516.4 STA_VDBB.scala 207:29:@15541.4 STA_VDBB.scala 207:29:@16308.4 STA_VDBB.scala 207:29:@16333.4 STA_VDBB.scala 207:29:@17100.4 STA_VDBB.scala 207:29:@17125.4 STA_VDBB.scala 207:29:@17892.4 STA_VDBB.scala 207:29:@17917.4 STA_VDBB.scala 207:29:@18684.4 STA_VDBB.scala 207:29:@18709.4 STA_VDBB.scala 241:23:@19019.4 STA_VDBB.scala 260:29:@19140.4 STA_VDBB.scala 260:29:@19165.4 STA_VDBB.scala 260:29:@19404.4 STA_VDBB.scala 260:29:@19429.4 STA_VDBB.scala 260:29:@19668.4 STA_VDBB.scala 260:29:@19693.4 STA_VDBB.scala 260:29:@19932.4 STA_VDBB.scala 260:29:@19957.4 STA_VDBB.scala 260:29:@20196.4 STA_VDBB.scala 260:29:@20221.4 STA_VDBB.scala 260:29:@20460.4 STA_VDBB.scala 260:29:@20485.4 STA_VDBB.scala 260:29:@20724.4 STA_VDBB.scala 260:29:@20749.4 STA_VDBB.scala 260:29:@20988.4 STA_VDBB.scala 260:29:@21013.4 STA_VDBB.scala 339:29:@21972.4 STA_VDBB.scala 339:29:@21997.4 STA_VDBB.scala 339:29:@22764.4 STA_VDBB.scala 339:29:@22789.4 STA_VDBB.scala 339:29:@23556.4 STA_VDBB.scala 339:29:@23581.4 STA_VDBB.scala 339:29:@24348.4 STA_VDBB.scala 339:29:@24373.4 STA_VDBB.scala 339:29:@25140.4 STA_VDBB.scala 339:29:@25165.4 STA_VDBB.scala 339:29:@25932.4 STA_VDBB.scala 339:29:@25957.4 STA_VDBB.scala 339:29:@26724.4 STA_VDBB.scala 339:29:@26749.4 STA_VDBB.scala 339:29:@27516.4 STA_VDBB.scala 339:29:@27541.4]
  assign ffb1_io_in_tag_1_0 = S8DP1_13_io_out_tag_0; // @[STA_VDBB.scala 108:23:@10204.4 STA_VDBB.scala 127:29:@10367.4 STA_VDBB.scala 127:29:@10392.4 STA_VDBB.scala 127:29:@10631.4 STA_VDBB.scala 127:29:@10656.4 STA_VDBB.scala 127:29:@10895.4 STA_VDBB.scala 127:29:@10920.4 STA_VDBB.scala 127:29:@11159.4 STA_VDBB.scala 127:29:@11184.4 STA_VDBB.scala 127:29:@11423.4 STA_VDBB.scala 127:29:@11448.4 STA_VDBB.scala 127:29:@11687.4 STA_VDBB.scala 127:29:@11712.4 STA_VDBB.scala 127:29:@11951.4 STA_VDBB.scala 127:29:@11976.4 STA_VDBB.scala 127:29:@12215.4 STA_VDBB.scala 127:29:@12240.4 STA_VDBB.scala 207:29:@13199.4 STA_VDBB.scala 207:29:@13224.4 STA_VDBB.scala 207:29:@13991.4 STA_VDBB.scala 207:29:@14016.4 STA_VDBB.scala 207:29:@14783.4 STA_VDBB.scala 207:29:@14808.4 STA_VDBB.scala 207:29:@15575.4 STA_VDBB.scala 207:29:@15600.4 STA_VDBB.scala 207:29:@16367.4 STA_VDBB.scala 207:29:@16392.4 STA_VDBB.scala 207:29:@17159.4 STA_VDBB.scala 207:29:@17184.4 STA_VDBB.scala 207:29:@17951.4 STA_VDBB.scala 207:29:@17976.4 STA_VDBB.scala 207:29:@18743.4 STA_VDBB.scala 207:29:@18768.4 STA_VDBB.scala 241:23:@19036.4 STA_VDBB.scala 260:29:@19199.4 STA_VDBB.scala 260:29:@19224.4 STA_VDBB.scala 260:29:@19463.4 STA_VDBB.scala 260:29:@19488.4 STA_VDBB.scala 260:29:@19727.4 STA_VDBB.scala 260:29:@19752.4 STA_VDBB.scala 260:29:@19991.4 STA_VDBB.scala 260:29:@20016.4 STA_VDBB.scala 260:29:@20255.4 STA_VDBB.scala 260:29:@20280.4 STA_VDBB.scala 260:29:@20519.4 STA_VDBB.scala 260:29:@20544.4 STA_VDBB.scala 260:29:@20783.4 STA_VDBB.scala 260:29:@20808.4 STA_VDBB.scala 260:29:@21047.4 STA_VDBB.scala 260:29:@21072.4 STA_VDBB.scala 339:29:@22031.4 STA_VDBB.scala 339:29:@22056.4 STA_VDBB.scala 339:29:@22823.4 STA_VDBB.scala 339:29:@22848.4 STA_VDBB.scala 339:29:@23615.4 STA_VDBB.scala 339:29:@23640.4 STA_VDBB.scala 339:29:@24407.4 STA_VDBB.scala 339:29:@24432.4 STA_VDBB.scala 339:29:@25199.4 STA_VDBB.scala 339:29:@25224.4 STA_VDBB.scala 339:29:@25991.4 STA_VDBB.scala 339:29:@26016.4 STA_VDBB.scala 339:29:@26783.4 STA_VDBB.scala 339:29:@26808.4 STA_VDBB.scala 339:29:@27575.4 STA_VDBB.scala 339:29:@27600.4]
  assign ffb1_io_in_tag_1_1 = S8DP1_13_io_out_tag_1; // @[STA_VDBB.scala 108:23:@10205.4 STA_VDBB.scala 127:29:@10368.4 STA_VDBB.scala 127:29:@10393.4 STA_VDBB.scala 127:29:@10632.4 STA_VDBB.scala 127:29:@10657.4 STA_VDBB.scala 127:29:@10896.4 STA_VDBB.scala 127:29:@10921.4 STA_VDBB.scala 127:29:@11160.4 STA_VDBB.scala 127:29:@11185.4 STA_VDBB.scala 127:29:@11424.4 STA_VDBB.scala 127:29:@11449.4 STA_VDBB.scala 127:29:@11688.4 STA_VDBB.scala 127:29:@11713.4 STA_VDBB.scala 127:29:@11952.4 STA_VDBB.scala 127:29:@11977.4 STA_VDBB.scala 127:29:@12216.4 STA_VDBB.scala 127:29:@12241.4 STA_VDBB.scala 207:29:@13200.4 STA_VDBB.scala 207:29:@13225.4 STA_VDBB.scala 207:29:@13992.4 STA_VDBB.scala 207:29:@14017.4 STA_VDBB.scala 207:29:@14784.4 STA_VDBB.scala 207:29:@14809.4 STA_VDBB.scala 207:29:@15576.4 STA_VDBB.scala 207:29:@15601.4 STA_VDBB.scala 207:29:@16368.4 STA_VDBB.scala 207:29:@16393.4 STA_VDBB.scala 207:29:@17160.4 STA_VDBB.scala 207:29:@17185.4 STA_VDBB.scala 207:29:@17952.4 STA_VDBB.scala 207:29:@17977.4 STA_VDBB.scala 207:29:@18744.4 STA_VDBB.scala 207:29:@18769.4 STA_VDBB.scala 241:23:@19037.4 STA_VDBB.scala 260:29:@19200.4 STA_VDBB.scala 260:29:@19225.4 STA_VDBB.scala 260:29:@19464.4 STA_VDBB.scala 260:29:@19489.4 STA_VDBB.scala 260:29:@19728.4 STA_VDBB.scala 260:29:@19753.4 STA_VDBB.scala 260:29:@19992.4 STA_VDBB.scala 260:29:@20017.4 STA_VDBB.scala 260:29:@20256.4 STA_VDBB.scala 260:29:@20281.4 STA_VDBB.scala 260:29:@20520.4 STA_VDBB.scala 260:29:@20545.4 STA_VDBB.scala 260:29:@20784.4 STA_VDBB.scala 260:29:@20809.4 STA_VDBB.scala 260:29:@21048.4 STA_VDBB.scala 260:29:@21073.4 STA_VDBB.scala 339:29:@22032.4 STA_VDBB.scala 339:29:@22057.4 STA_VDBB.scala 339:29:@22824.4 STA_VDBB.scala 339:29:@22849.4 STA_VDBB.scala 339:29:@23616.4 STA_VDBB.scala 339:29:@23641.4 STA_VDBB.scala 339:29:@24408.4 STA_VDBB.scala 339:29:@24433.4 STA_VDBB.scala 339:29:@25200.4 STA_VDBB.scala 339:29:@25225.4 STA_VDBB.scala 339:29:@25992.4 STA_VDBB.scala 339:29:@26017.4 STA_VDBB.scala 339:29:@26784.4 STA_VDBB.scala 339:29:@26809.4 STA_VDBB.scala 339:29:@27576.4 STA_VDBB.scala 339:29:@27601.4]
  assign ffb1_io_in_tag_1_2 = S8DP1_13_io_out_tag_2; // @[STA_VDBB.scala 108:23:@10206.4 STA_VDBB.scala 127:29:@10369.4 STA_VDBB.scala 127:29:@10394.4 STA_VDBB.scala 127:29:@10633.4 STA_VDBB.scala 127:29:@10658.4 STA_VDBB.scala 127:29:@10897.4 STA_VDBB.scala 127:29:@10922.4 STA_VDBB.scala 127:29:@11161.4 STA_VDBB.scala 127:29:@11186.4 STA_VDBB.scala 127:29:@11425.4 STA_VDBB.scala 127:29:@11450.4 STA_VDBB.scala 127:29:@11689.4 STA_VDBB.scala 127:29:@11714.4 STA_VDBB.scala 127:29:@11953.4 STA_VDBB.scala 127:29:@11978.4 STA_VDBB.scala 127:29:@12217.4 STA_VDBB.scala 127:29:@12242.4 STA_VDBB.scala 207:29:@13201.4 STA_VDBB.scala 207:29:@13226.4 STA_VDBB.scala 207:29:@13993.4 STA_VDBB.scala 207:29:@14018.4 STA_VDBB.scala 207:29:@14785.4 STA_VDBB.scala 207:29:@14810.4 STA_VDBB.scala 207:29:@15577.4 STA_VDBB.scala 207:29:@15602.4 STA_VDBB.scala 207:29:@16369.4 STA_VDBB.scala 207:29:@16394.4 STA_VDBB.scala 207:29:@17161.4 STA_VDBB.scala 207:29:@17186.4 STA_VDBB.scala 207:29:@17953.4 STA_VDBB.scala 207:29:@17978.4 STA_VDBB.scala 207:29:@18745.4 STA_VDBB.scala 207:29:@18770.4 STA_VDBB.scala 241:23:@19038.4 STA_VDBB.scala 260:29:@19201.4 STA_VDBB.scala 260:29:@19226.4 STA_VDBB.scala 260:29:@19465.4 STA_VDBB.scala 260:29:@19490.4 STA_VDBB.scala 260:29:@19729.4 STA_VDBB.scala 260:29:@19754.4 STA_VDBB.scala 260:29:@19993.4 STA_VDBB.scala 260:29:@20018.4 STA_VDBB.scala 260:29:@20257.4 STA_VDBB.scala 260:29:@20282.4 STA_VDBB.scala 260:29:@20521.4 STA_VDBB.scala 260:29:@20546.4 STA_VDBB.scala 260:29:@20785.4 STA_VDBB.scala 260:29:@20810.4 STA_VDBB.scala 260:29:@21049.4 STA_VDBB.scala 260:29:@21074.4 STA_VDBB.scala 339:29:@22033.4 STA_VDBB.scala 339:29:@22058.4 STA_VDBB.scala 339:29:@22825.4 STA_VDBB.scala 339:29:@22850.4 STA_VDBB.scala 339:29:@23617.4 STA_VDBB.scala 339:29:@23642.4 STA_VDBB.scala 339:29:@24409.4 STA_VDBB.scala 339:29:@24434.4 STA_VDBB.scala 339:29:@25201.4 STA_VDBB.scala 339:29:@25226.4 STA_VDBB.scala 339:29:@25993.4 STA_VDBB.scala 339:29:@26018.4 STA_VDBB.scala 339:29:@26785.4 STA_VDBB.scala 339:29:@26810.4 STA_VDBB.scala 339:29:@27577.4 STA_VDBB.scala 339:29:@27602.4]
  assign ffb1_io_in_tag_1_3 = S8DP1_13_io_out_tag_3; // @[STA_VDBB.scala 108:23:@10207.4 STA_VDBB.scala 127:29:@10370.4 STA_VDBB.scala 127:29:@10395.4 STA_VDBB.scala 127:29:@10634.4 STA_VDBB.scala 127:29:@10659.4 STA_VDBB.scala 127:29:@10898.4 STA_VDBB.scala 127:29:@10923.4 STA_VDBB.scala 127:29:@11162.4 STA_VDBB.scala 127:29:@11187.4 STA_VDBB.scala 127:29:@11426.4 STA_VDBB.scala 127:29:@11451.4 STA_VDBB.scala 127:29:@11690.4 STA_VDBB.scala 127:29:@11715.4 STA_VDBB.scala 127:29:@11954.4 STA_VDBB.scala 127:29:@11979.4 STA_VDBB.scala 127:29:@12218.4 STA_VDBB.scala 127:29:@12243.4 STA_VDBB.scala 207:29:@13202.4 STA_VDBB.scala 207:29:@13227.4 STA_VDBB.scala 207:29:@13994.4 STA_VDBB.scala 207:29:@14019.4 STA_VDBB.scala 207:29:@14786.4 STA_VDBB.scala 207:29:@14811.4 STA_VDBB.scala 207:29:@15578.4 STA_VDBB.scala 207:29:@15603.4 STA_VDBB.scala 207:29:@16370.4 STA_VDBB.scala 207:29:@16395.4 STA_VDBB.scala 207:29:@17162.4 STA_VDBB.scala 207:29:@17187.4 STA_VDBB.scala 207:29:@17954.4 STA_VDBB.scala 207:29:@17979.4 STA_VDBB.scala 207:29:@18746.4 STA_VDBB.scala 207:29:@18771.4 STA_VDBB.scala 241:23:@19039.4 STA_VDBB.scala 260:29:@19202.4 STA_VDBB.scala 260:29:@19227.4 STA_VDBB.scala 260:29:@19466.4 STA_VDBB.scala 260:29:@19491.4 STA_VDBB.scala 260:29:@19730.4 STA_VDBB.scala 260:29:@19755.4 STA_VDBB.scala 260:29:@19994.4 STA_VDBB.scala 260:29:@20019.4 STA_VDBB.scala 260:29:@20258.4 STA_VDBB.scala 260:29:@20283.4 STA_VDBB.scala 260:29:@20522.4 STA_VDBB.scala 260:29:@20547.4 STA_VDBB.scala 260:29:@20786.4 STA_VDBB.scala 260:29:@20811.4 STA_VDBB.scala 260:29:@21050.4 STA_VDBB.scala 260:29:@21075.4 STA_VDBB.scala 339:29:@22034.4 STA_VDBB.scala 339:29:@22059.4 STA_VDBB.scala 339:29:@22826.4 STA_VDBB.scala 339:29:@22851.4 STA_VDBB.scala 339:29:@23618.4 STA_VDBB.scala 339:29:@23643.4 STA_VDBB.scala 339:29:@24410.4 STA_VDBB.scala 339:29:@24435.4 STA_VDBB.scala 339:29:@25202.4 STA_VDBB.scala 339:29:@25227.4 STA_VDBB.scala 339:29:@25994.4 STA_VDBB.scala 339:29:@26019.4 STA_VDBB.scala 339:29:@26786.4 STA_VDBB.scala 339:29:@26811.4 STA_VDBB.scala 339:29:@27578.4 STA_VDBB.scala 339:29:@27603.4]
  assign ffb1_io_in_tag_1_4 = S8DP1_13_io_out_tag_4; // @[STA_VDBB.scala 108:23:@10208.4 STA_VDBB.scala 127:29:@10371.4 STA_VDBB.scala 127:29:@10396.4 STA_VDBB.scala 127:29:@10635.4 STA_VDBB.scala 127:29:@10660.4 STA_VDBB.scala 127:29:@10899.4 STA_VDBB.scala 127:29:@10924.4 STA_VDBB.scala 127:29:@11163.4 STA_VDBB.scala 127:29:@11188.4 STA_VDBB.scala 127:29:@11427.4 STA_VDBB.scala 127:29:@11452.4 STA_VDBB.scala 127:29:@11691.4 STA_VDBB.scala 127:29:@11716.4 STA_VDBB.scala 127:29:@11955.4 STA_VDBB.scala 127:29:@11980.4 STA_VDBB.scala 127:29:@12219.4 STA_VDBB.scala 127:29:@12244.4 STA_VDBB.scala 207:29:@13203.4 STA_VDBB.scala 207:29:@13228.4 STA_VDBB.scala 207:29:@13995.4 STA_VDBB.scala 207:29:@14020.4 STA_VDBB.scala 207:29:@14787.4 STA_VDBB.scala 207:29:@14812.4 STA_VDBB.scala 207:29:@15579.4 STA_VDBB.scala 207:29:@15604.4 STA_VDBB.scala 207:29:@16371.4 STA_VDBB.scala 207:29:@16396.4 STA_VDBB.scala 207:29:@17163.4 STA_VDBB.scala 207:29:@17188.4 STA_VDBB.scala 207:29:@17955.4 STA_VDBB.scala 207:29:@17980.4 STA_VDBB.scala 207:29:@18747.4 STA_VDBB.scala 207:29:@18772.4 STA_VDBB.scala 241:23:@19040.4 STA_VDBB.scala 260:29:@19203.4 STA_VDBB.scala 260:29:@19228.4 STA_VDBB.scala 260:29:@19467.4 STA_VDBB.scala 260:29:@19492.4 STA_VDBB.scala 260:29:@19731.4 STA_VDBB.scala 260:29:@19756.4 STA_VDBB.scala 260:29:@19995.4 STA_VDBB.scala 260:29:@20020.4 STA_VDBB.scala 260:29:@20259.4 STA_VDBB.scala 260:29:@20284.4 STA_VDBB.scala 260:29:@20523.4 STA_VDBB.scala 260:29:@20548.4 STA_VDBB.scala 260:29:@20787.4 STA_VDBB.scala 260:29:@20812.4 STA_VDBB.scala 260:29:@21051.4 STA_VDBB.scala 260:29:@21076.4 STA_VDBB.scala 339:29:@22035.4 STA_VDBB.scala 339:29:@22060.4 STA_VDBB.scala 339:29:@22827.4 STA_VDBB.scala 339:29:@22852.4 STA_VDBB.scala 339:29:@23619.4 STA_VDBB.scala 339:29:@23644.4 STA_VDBB.scala 339:29:@24411.4 STA_VDBB.scala 339:29:@24436.4 STA_VDBB.scala 339:29:@25203.4 STA_VDBB.scala 339:29:@25228.4 STA_VDBB.scala 339:29:@25995.4 STA_VDBB.scala 339:29:@26020.4 STA_VDBB.scala 339:29:@26787.4 STA_VDBB.scala 339:29:@26812.4 STA_VDBB.scala 339:29:@27579.4 STA_VDBB.scala 339:29:@27604.4]
  assign ffb1_io_in_tag_1_5 = S8DP1_13_io_out_tag_5; // @[STA_VDBB.scala 108:23:@10209.4 STA_VDBB.scala 127:29:@10372.4 STA_VDBB.scala 127:29:@10397.4 STA_VDBB.scala 127:29:@10636.4 STA_VDBB.scala 127:29:@10661.4 STA_VDBB.scala 127:29:@10900.4 STA_VDBB.scala 127:29:@10925.4 STA_VDBB.scala 127:29:@11164.4 STA_VDBB.scala 127:29:@11189.4 STA_VDBB.scala 127:29:@11428.4 STA_VDBB.scala 127:29:@11453.4 STA_VDBB.scala 127:29:@11692.4 STA_VDBB.scala 127:29:@11717.4 STA_VDBB.scala 127:29:@11956.4 STA_VDBB.scala 127:29:@11981.4 STA_VDBB.scala 127:29:@12220.4 STA_VDBB.scala 127:29:@12245.4 STA_VDBB.scala 207:29:@13204.4 STA_VDBB.scala 207:29:@13229.4 STA_VDBB.scala 207:29:@13996.4 STA_VDBB.scala 207:29:@14021.4 STA_VDBB.scala 207:29:@14788.4 STA_VDBB.scala 207:29:@14813.4 STA_VDBB.scala 207:29:@15580.4 STA_VDBB.scala 207:29:@15605.4 STA_VDBB.scala 207:29:@16372.4 STA_VDBB.scala 207:29:@16397.4 STA_VDBB.scala 207:29:@17164.4 STA_VDBB.scala 207:29:@17189.4 STA_VDBB.scala 207:29:@17956.4 STA_VDBB.scala 207:29:@17981.4 STA_VDBB.scala 207:29:@18748.4 STA_VDBB.scala 207:29:@18773.4 STA_VDBB.scala 241:23:@19041.4 STA_VDBB.scala 260:29:@19204.4 STA_VDBB.scala 260:29:@19229.4 STA_VDBB.scala 260:29:@19468.4 STA_VDBB.scala 260:29:@19493.4 STA_VDBB.scala 260:29:@19732.4 STA_VDBB.scala 260:29:@19757.4 STA_VDBB.scala 260:29:@19996.4 STA_VDBB.scala 260:29:@20021.4 STA_VDBB.scala 260:29:@20260.4 STA_VDBB.scala 260:29:@20285.4 STA_VDBB.scala 260:29:@20524.4 STA_VDBB.scala 260:29:@20549.4 STA_VDBB.scala 260:29:@20788.4 STA_VDBB.scala 260:29:@20813.4 STA_VDBB.scala 260:29:@21052.4 STA_VDBB.scala 260:29:@21077.4 STA_VDBB.scala 339:29:@22036.4 STA_VDBB.scala 339:29:@22061.4 STA_VDBB.scala 339:29:@22828.4 STA_VDBB.scala 339:29:@22853.4 STA_VDBB.scala 339:29:@23620.4 STA_VDBB.scala 339:29:@23645.4 STA_VDBB.scala 339:29:@24412.4 STA_VDBB.scala 339:29:@24437.4 STA_VDBB.scala 339:29:@25204.4 STA_VDBB.scala 339:29:@25229.4 STA_VDBB.scala 339:29:@25996.4 STA_VDBB.scala 339:29:@26021.4 STA_VDBB.scala 339:29:@26788.4 STA_VDBB.scala 339:29:@26813.4 STA_VDBB.scala 339:29:@27580.4 STA_VDBB.scala 339:29:@27605.4]
  assign ffb1_io_in_tag_1_6 = S8DP1_13_io_out_tag_6; // @[STA_VDBB.scala 108:23:@10210.4 STA_VDBB.scala 127:29:@10373.4 STA_VDBB.scala 127:29:@10398.4 STA_VDBB.scala 127:29:@10637.4 STA_VDBB.scala 127:29:@10662.4 STA_VDBB.scala 127:29:@10901.4 STA_VDBB.scala 127:29:@10926.4 STA_VDBB.scala 127:29:@11165.4 STA_VDBB.scala 127:29:@11190.4 STA_VDBB.scala 127:29:@11429.4 STA_VDBB.scala 127:29:@11454.4 STA_VDBB.scala 127:29:@11693.4 STA_VDBB.scala 127:29:@11718.4 STA_VDBB.scala 127:29:@11957.4 STA_VDBB.scala 127:29:@11982.4 STA_VDBB.scala 127:29:@12221.4 STA_VDBB.scala 127:29:@12246.4 STA_VDBB.scala 207:29:@13205.4 STA_VDBB.scala 207:29:@13230.4 STA_VDBB.scala 207:29:@13997.4 STA_VDBB.scala 207:29:@14022.4 STA_VDBB.scala 207:29:@14789.4 STA_VDBB.scala 207:29:@14814.4 STA_VDBB.scala 207:29:@15581.4 STA_VDBB.scala 207:29:@15606.4 STA_VDBB.scala 207:29:@16373.4 STA_VDBB.scala 207:29:@16398.4 STA_VDBB.scala 207:29:@17165.4 STA_VDBB.scala 207:29:@17190.4 STA_VDBB.scala 207:29:@17957.4 STA_VDBB.scala 207:29:@17982.4 STA_VDBB.scala 207:29:@18749.4 STA_VDBB.scala 207:29:@18774.4 STA_VDBB.scala 241:23:@19042.4 STA_VDBB.scala 260:29:@19205.4 STA_VDBB.scala 260:29:@19230.4 STA_VDBB.scala 260:29:@19469.4 STA_VDBB.scala 260:29:@19494.4 STA_VDBB.scala 260:29:@19733.4 STA_VDBB.scala 260:29:@19758.4 STA_VDBB.scala 260:29:@19997.4 STA_VDBB.scala 260:29:@20022.4 STA_VDBB.scala 260:29:@20261.4 STA_VDBB.scala 260:29:@20286.4 STA_VDBB.scala 260:29:@20525.4 STA_VDBB.scala 260:29:@20550.4 STA_VDBB.scala 260:29:@20789.4 STA_VDBB.scala 260:29:@20814.4 STA_VDBB.scala 260:29:@21053.4 STA_VDBB.scala 260:29:@21078.4 STA_VDBB.scala 339:29:@22037.4 STA_VDBB.scala 339:29:@22062.4 STA_VDBB.scala 339:29:@22829.4 STA_VDBB.scala 339:29:@22854.4 STA_VDBB.scala 339:29:@23621.4 STA_VDBB.scala 339:29:@23646.4 STA_VDBB.scala 339:29:@24413.4 STA_VDBB.scala 339:29:@24438.4 STA_VDBB.scala 339:29:@25205.4 STA_VDBB.scala 339:29:@25230.4 STA_VDBB.scala 339:29:@25997.4 STA_VDBB.scala 339:29:@26022.4 STA_VDBB.scala 339:29:@26789.4 STA_VDBB.scala 339:29:@26814.4 STA_VDBB.scala 339:29:@27581.4 STA_VDBB.scala 339:29:@27606.4]
  assign ffb1_io_in_tag_1_7 = S8DP1_13_io_out_tag_7; // @[STA_VDBB.scala 108:23:@10211.4 STA_VDBB.scala 127:29:@10374.4 STA_VDBB.scala 127:29:@10399.4 STA_VDBB.scala 127:29:@10638.4 STA_VDBB.scala 127:29:@10663.4 STA_VDBB.scala 127:29:@10902.4 STA_VDBB.scala 127:29:@10927.4 STA_VDBB.scala 127:29:@11166.4 STA_VDBB.scala 127:29:@11191.4 STA_VDBB.scala 127:29:@11430.4 STA_VDBB.scala 127:29:@11455.4 STA_VDBB.scala 127:29:@11694.4 STA_VDBB.scala 127:29:@11719.4 STA_VDBB.scala 127:29:@11958.4 STA_VDBB.scala 127:29:@11983.4 STA_VDBB.scala 127:29:@12222.4 STA_VDBB.scala 127:29:@12247.4 STA_VDBB.scala 207:29:@13206.4 STA_VDBB.scala 207:29:@13231.4 STA_VDBB.scala 207:29:@13998.4 STA_VDBB.scala 207:29:@14023.4 STA_VDBB.scala 207:29:@14790.4 STA_VDBB.scala 207:29:@14815.4 STA_VDBB.scala 207:29:@15582.4 STA_VDBB.scala 207:29:@15607.4 STA_VDBB.scala 207:29:@16374.4 STA_VDBB.scala 207:29:@16399.4 STA_VDBB.scala 207:29:@17166.4 STA_VDBB.scala 207:29:@17191.4 STA_VDBB.scala 207:29:@17958.4 STA_VDBB.scala 207:29:@17983.4 STA_VDBB.scala 207:29:@18750.4 STA_VDBB.scala 207:29:@18775.4 STA_VDBB.scala 241:23:@19043.4 STA_VDBB.scala 260:29:@19206.4 STA_VDBB.scala 260:29:@19231.4 STA_VDBB.scala 260:29:@19470.4 STA_VDBB.scala 260:29:@19495.4 STA_VDBB.scala 260:29:@19734.4 STA_VDBB.scala 260:29:@19759.4 STA_VDBB.scala 260:29:@19998.4 STA_VDBB.scala 260:29:@20023.4 STA_VDBB.scala 260:29:@20262.4 STA_VDBB.scala 260:29:@20287.4 STA_VDBB.scala 260:29:@20526.4 STA_VDBB.scala 260:29:@20551.4 STA_VDBB.scala 260:29:@20790.4 STA_VDBB.scala 260:29:@20815.4 STA_VDBB.scala 260:29:@21054.4 STA_VDBB.scala 260:29:@21079.4 STA_VDBB.scala 339:29:@22038.4 STA_VDBB.scala 339:29:@22063.4 STA_VDBB.scala 339:29:@22830.4 STA_VDBB.scala 339:29:@22855.4 STA_VDBB.scala 339:29:@23622.4 STA_VDBB.scala 339:29:@23647.4 STA_VDBB.scala 339:29:@24414.4 STA_VDBB.scala 339:29:@24439.4 STA_VDBB.scala 339:29:@25206.4 STA_VDBB.scala 339:29:@25231.4 STA_VDBB.scala 339:29:@25998.4 STA_VDBB.scala 339:29:@26023.4 STA_VDBB.scala 339:29:@26790.4 STA_VDBB.scala 339:29:@26815.4 STA_VDBB.scala 339:29:@27582.4 STA_VDBB.scala 339:29:@27607.4]
  assign ffb1_io_in_tag_2_0 = S8DP1_14_io_out_tag_0; // @[STA_VDBB.scala 108:23:@10228.4 STA_VDBB.scala 127:29:@10433.4 STA_VDBB.scala 127:29:@10458.4 STA_VDBB.scala 127:29:@10697.4 STA_VDBB.scala 127:29:@10722.4 STA_VDBB.scala 127:29:@10961.4 STA_VDBB.scala 127:29:@10986.4 STA_VDBB.scala 127:29:@11225.4 STA_VDBB.scala 127:29:@11250.4 STA_VDBB.scala 127:29:@11489.4 STA_VDBB.scala 127:29:@11514.4 STA_VDBB.scala 127:29:@11753.4 STA_VDBB.scala 127:29:@11778.4 STA_VDBB.scala 127:29:@12017.4 STA_VDBB.scala 127:29:@12042.4 STA_VDBB.scala 127:29:@12281.4 STA_VDBB.scala 127:29:@12306.4 STA_VDBB.scala 207:29:@13265.4 STA_VDBB.scala 207:29:@13290.4 STA_VDBB.scala 207:29:@14057.4 STA_VDBB.scala 207:29:@14082.4 STA_VDBB.scala 207:29:@14849.4 STA_VDBB.scala 207:29:@14874.4 STA_VDBB.scala 207:29:@15641.4 STA_VDBB.scala 207:29:@15666.4 STA_VDBB.scala 207:29:@16433.4 STA_VDBB.scala 207:29:@16458.4 STA_VDBB.scala 207:29:@17225.4 STA_VDBB.scala 207:29:@17250.4 STA_VDBB.scala 207:29:@18017.4 STA_VDBB.scala 207:29:@18042.4 STA_VDBB.scala 207:29:@18809.4 STA_VDBB.scala 207:29:@18834.4 STA_VDBB.scala 241:23:@19060.4 STA_VDBB.scala 260:29:@19265.4 STA_VDBB.scala 260:29:@19290.4 STA_VDBB.scala 260:29:@19529.4 STA_VDBB.scala 260:29:@19554.4 STA_VDBB.scala 260:29:@19793.4 STA_VDBB.scala 260:29:@19818.4 STA_VDBB.scala 260:29:@20057.4 STA_VDBB.scala 260:29:@20082.4 STA_VDBB.scala 260:29:@20321.4 STA_VDBB.scala 260:29:@20346.4 STA_VDBB.scala 260:29:@20585.4 STA_VDBB.scala 260:29:@20610.4 STA_VDBB.scala 260:29:@20849.4 STA_VDBB.scala 260:29:@20874.4 STA_VDBB.scala 260:29:@21113.4 STA_VDBB.scala 260:29:@21138.4 STA_VDBB.scala 339:29:@22097.4 STA_VDBB.scala 339:29:@22122.4 STA_VDBB.scala 339:29:@22889.4 STA_VDBB.scala 339:29:@22914.4 STA_VDBB.scala 339:29:@23681.4 STA_VDBB.scala 339:29:@23706.4 STA_VDBB.scala 339:29:@24473.4 STA_VDBB.scala 339:29:@24498.4 STA_VDBB.scala 339:29:@25265.4 STA_VDBB.scala 339:29:@25290.4 STA_VDBB.scala 339:29:@26057.4 STA_VDBB.scala 339:29:@26082.4 STA_VDBB.scala 339:29:@26849.4 STA_VDBB.scala 339:29:@26874.4 STA_VDBB.scala 339:29:@27641.4 STA_VDBB.scala 339:29:@27666.4]
  assign ffb1_io_in_tag_2_1 = S8DP1_14_io_out_tag_1; // @[STA_VDBB.scala 108:23:@10229.4 STA_VDBB.scala 127:29:@10434.4 STA_VDBB.scala 127:29:@10459.4 STA_VDBB.scala 127:29:@10698.4 STA_VDBB.scala 127:29:@10723.4 STA_VDBB.scala 127:29:@10962.4 STA_VDBB.scala 127:29:@10987.4 STA_VDBB.scala 127:29:@11226.4 STA_VDBB.scala 127:29:@11251.4 STA_VDBB.scala 127:29:@11490.4 STA_VDBB.scala 127:29:@11515.4 STA_VDBB.scala 127:29:@11754.4 STA_VDBB.scala 127:29:@11779.4 STA_VDBB.scala 127:29:@12018.4 STA_VDBB.scala 127:29:@12043.4 STA_VDBB.scala 127:29:@12282.4 STA_VDBB.scala 127:29:@12307.4 STA_VDBB.scala 207:29:@13266.4 STA_VDBB.scala 207:29:@13291.4 STA_VDBB.scala 207:29:@14058.4 STA_VDBB.scala 207:29:@14083.4 STA_VDBB.scala 207:29:@14850.4 STA_VDBB.scala 207:29:@14875.4 STA_VDBB.scala 207:29:@15642.4 STA_VDBB.scala 207:29:@15667.4 STA_VDBB.scala 207:29:@16434.4 STA_VDBB.scala 207:29:@16459.4 STA_VDBB.scala 207:29:@17226.4 STA_VDBB.scala 207:29:@17251.4 STA_VDBB.scala 207:29:@18018.4 STA_VDBB.scala 207:29:@18043.4 STA_VDBB.scala 207:29:@18810.4 STA_VDBB.scala 207:29:@18835.4 STA_VDBB.scala 241:23:@19061.4 STA_VDBB.scala 260:29:@19266.4 STA_VDBB.scala 260:29:@19291.4 STA_VDBB.scala 260:29:@19530.4 STA_VDBB.scala 260:29:@19555.4 STA_VDBB.scala 260:29:@19794.4 STA_VDBB.scala 260:29:@19819.4 STA_VDBB.scala 260:29:@20058.4 STA_VDBB.scala 260:29:@20083.4 STA_VDBB.scala 260:29:@20322.4 STA_VDBB.scala 260:29:@20347.4 STA_VDBB.scala 260:29:@20586.4 STA_VDBB.scala 260:29:@20611.4 STA_VDBB.scala 260:29:@20850.4 STA_VDBB.scala 260:29:@20875.4 STA_VDBB.scala 260:29:@21114.4 STA_VDBB.scala 260:29:@21139.4 STA_VDBB.scala 339:29:@22098.4 STA_VDBB.scala 339:29:@22123.4 STA_VDBB.scala 339:29:@22890.4 STA_VDBB.scala 339:29:@22915.4 STA_VDBB.scala 339:29:@23682.4 STA_VDBB.scala 339:29:@23707.4 STA_VDBB.scala 339:29:@24474.4 STA_VDBB.scala 339:29:@24499.4 STA_VDBB.scala 339:29:@25266.4 STA_VDBB.scala 339:29:@25291.4 STA_VDBB.scala 339:29:@26058.4 STA_VDBB.scala 339:29:@26083.4 STA_VDBB.scala 339:29:@26850.4 STA_VDBB.scala 339:29:@26875.4 STA_VDBB.scala 339:29:@27642.4 STA_VDBB.scala 339:29:@27667.4]
  assign ffb1_io_in_tag_2_2 = S8DP1_14_io_out_tag_2; // @[STA_VDBB.scala 108:23:@10230.4 STA_VDBB.scala 127:29:@10435.4 STA_VDBB.scala 127:29:@10460.4 STA_VDBB.scala 127:29:@10699.4 STA_VDBB.scala 127:29:@10724.4 STA_VDBB.scala 127:29:@10963.4 STA_VDBB.scala 127:29:@10988.4 STA_VDBB.scala 127:29:@11227.4 STA_VDBB.scala 127:29:@11252.4 STA_VDBB.scala 127:29:@11491.4 STA_VDBB.scala 127:29:@11516.4 STA_VDBB.scala 127:29:@11755.4 STA_VDBB.scala 127:29:@11780.4 STA_VDBB.scala 127:29:@12019.4 STA_VDBB.scala 127:29:@12044.4 STA_VDBB.scala 127:29:@12283.4 STA_VDBB.scala 127:29:@12308.4 STA_VDBB.scala 207:29:@13267.4 STA_VDBB.scala 207:29:@13292.4 STA_VDBB.scala 207:29:@14059.4 STA_VDBB.scala 207:29:@14084.4 STA_VDBB.scala 207:29:@14851.4 STA_VDBB.scala 207:29:@14876.4 STA_VDBB.scala 207:29:@15643.4 STA_VDBB.scala 207:29:@15668.4 STA_VDBB.scala 207:29:@16435.4 STA_VDBB.scala 207:29:@16460.4 STA_VDBB.scala 207:29:@17227.4 STA_VDBB.scala 207:29:@17252.4 STA_VDBB.scala 207:29:@18019.4 STA_VDBB.scala 207:29:@18044.4 STA_VDBB.scala 207:29:@18811.4 STA_VDBB.scala 207:29:@18836.4 STA_VDBB.scala 241:23:@19062.4 STA_VDBB.scala 260:29:@19267.4 STA_VDBB.scala 260:29:@19292.4 STA_VDBB.scala 260:29:@19531.4 STA_VDBB.scala 260:29:@19556.4 STA_VDBB.scala 260:29:@19795.4 STA_VDBB.scala 260:29:@19820.4 STA_VDBB.scala 260:29:@20059.4 STA_VDBB.scala 260:29:@20084.4 STA_VDBB.scala 260:29:@20323.4 STA_VDBB.scala 260:29:@20348.4 STA_VDBB.scala 260:29:@20587.4 STA_VDBB.scala 260:29:@20612.4 STA_VDBB.scala 260:29:@20851.4 STA_VDBB.scala 260:29:@20876.4 STA_VDBB.scala 260:29:@21115.4 STA_VDBB.scala 260:29:@21140.4 STA_VDBB.scala 339:29:@22099.4 STA_VDBB.scala 339:29:@22124.4 STA_VDBB.scala 339:29:@22891.4 STA_VDBB.scala 339:29:@22916.4 STA_VDBB.scala 339:29:@23683.4 STA_VDBB.scala 339:29:@23708.4 STA_VDBB.scala 339:29:@24475.4 STA_VDBB.scala 339:29:@24500.4 STA_VDBB.scala 339:29:@25267.4 STA_VDBB.scala 339:29:@25292.4 STA_VDBB.scala 339:29:@26059.4 STA_VDBB.scala 339:29:@26084.4 STA_VDBB.scala 339:29:@26851.4 STA_VDBB.scala 339:29:@26876.4 STA_VDBB.scala 339:29:@27643.4 STA_VDBB.scala 339:29:@27668.4]
  assign ffb1_io_in_tag_2_3 = S8DP1_14_io_out_tag_3; // @[STA_VDBB.scala 108:23:@10231.4 STA_VDBB.scala 127:29:@10436.4 STA_VDBB.scala 127:29:@10461.4 STA_VDBB.scala 127:29:@10700.4 STA_VDBB.scala 127:29:@10725.4 STA_VDBB.scala 127:29:@10964.4 STA_VDBB.scala 127:29:@10989.4 STA_VDBB.scala 127:29:@11228.4 STA_VDBB.scala 127:29:@11253.4 STA_VDBB.scala 127:29:@11492.4 STA_VDBB.scala 127:29:@11517.4 STA_VDBB.scala 127:29:@11756.4 STA_VDBB.scala 127:29:@11781.4 STA_VDBB.scala 127:29:@12020.4 STA_VDBB.scala 127:29:@12045.4 STA_VDBB.scala 127:29:@12284.4 STA_VDBB.scala 127:29:@12309.4 STA_VDBB.scala 207:29:@13268.4 STA_VDBB.scala 207:29:@13293.4 STA_VDBB.scala 207:29:@14060.4 STA_VDBB.scala 207:29:@14085.4 STA_VDBB.scala 207:29:@14852.4 STA_VDBB.scala 207:29:@14877.4 STA_VDBB.scala 207:29:@15644.4 STA_VDBB.scala 207:29:@15669.4 STA_VDBB.scala 207:29:@16436.4 STA_VDBB.scala 207:29:@16461.4 STA_VDBB.scala 207:29:@17228.4 STA_VDBB.scala 207:29:@17253.4 STA_VDBB.scala 207:29:@18020.4 STA_VDBB.scala 207:29:@18045.4 STA_VDBB.scala 207:29:@18812.4 STA_VDBB.scala 207:29:@18837.4 STA_VDBB.scala 241:23:@19063.4 STA_VDBB.scala 260:29:@19268.4 STA_VDBB.scala 260:29:@19293.4 STA_VDBB.scala 260:29:@19532.4 STA_VDBB.scala 260:29:@19557.4 STA_VDBB.scala 260:29:@19796.4 STA_VDBB.scala 260:29:@19821.4 STA_VDBB.scala 260:29:@20060.4 STA_VDBB.scala 260:29:@20085.4 STA_VDBB.scala 260:29:@20324.4 STA_VDBB.scala 260:29:@20349.4 STA_VDBB.scala 260:29:@20588.4 STA_VDBB.scala 260:29:@20613.4 STA_VDBB.scala 260:29:@20852.4 STA_VDBB.scala 260:29:@20877.4 STA_VDBB.scala 260:29:@21116.4 STA_VDBB.scala 260:29:@21141.4 STA_VDBB.scala 339:29:@22100.4 STA_VDBB.scala 339:29:@22125.4 STA_VDBB.scala 339:29:@22892.4 STA_VDBB.scala 339:29:@22917.4 STA_VDBB.scala 339:29:@23684.4 STA_VDBB.scala 339:29:@23709.4 STA_VDBB.scala 339:29:@24476.4 STA_VDBB.scala 339:29:@24501.4 STA_VDBB.scala 339:29:@25268.4 STA_VDBB.scala 339:29:@25293.4 STA_VDBB.scala 339:29:@26060.4 STA_VDBB.scala 339:29:@26085.4 STA_VDBB.scala 339:29:@26852.4 STA_VDBB.scala 339:29:@26877.4 STA_VDBB.scala 339:29:@27644.4 STA_VDBB.scala 339:29:@27669.4]
  assign ffb1_io_in_tag_2_4 = S8DP1_14_io_out_tag_4; // @[STA_VDBB.scala 108:23:@10232.4 STA_VDBB.scala 127:29:@10437.4 STA_VDBB.scala 127:29:@10462.4 STA_VDBB.scala 127:29:@10701.4 STA_VDBB.scala 127:29:@10726.4 STA_VDBB.scala 127:29:@10965.4 STA_VDBB.scala 127:29:@10990.4 STA_VDBB.scala 127:29:@11229.4 STA_VDBB.scala 127:29:@11254.4 STA_VDBB.scala 127:29:@11493.4 STA_VDBB.scala 127:29:@11518.4 STA_VDBB.scala 127:29:@11757.4 STA_VDBB.scala 127:29:@11782.4 STA_VDBB.scala 127:29:@12021.4 STA_VDBB.scala 127:29:@12046.4 STA_VDBB.scala 127:29:@12285.4 STA_VDBB.scala 127:29:@12310.4 STA_VDBB.scala 207:29:@13269.4 STA_VDBB.scala 207:29:@13294.4 STA_VDBB.scala 207:29:@14061.4 STA_VDBB.scala 207:29:@14086.4 STA_VDBB.scala 207:29:@14853.4 STA_VDBB.scala 207:29:@14878.4 STA_VDBB.scala 207:29:@15645.4 STA_VDBB.scala 207:29:@15670.4 STA_VDBB.scala 207:29:@16437.4 STA_VDBB.scala 207:29:@16462.4 STA_VDBB.scala 207:29:@17229.4 STA_VDBB.scala 207:29:@17254.4 STA_VDBB.scala 207:29:@18021.4 STA_VDBB.scala 207:29:@18046.4 STA_VDBB.scala 207:29:@18813.4 STA_VDBB.scala 207:29:@18838.4 STA_VDBB.scala 241:23:@19064.4 STA_VDBB.scala 260:29:@19269.4 STA_VDBB.scala 260:29:@19294.4 STA_VDBB.scala 260:29:@19533.4 STA_VDBB.scala 260:29:@19558.4 STA_VDBB.scala 260:29:@19797.4 STA_VDBB.scala 260:29:@19822.4 STA_VDBB.scala 260:29:@20061.4 STA_VDBB.scala 260:29:@20086.4 STA_VDBB.scala 260:29:@20325.4 STA_VDBB.scala 260:29:@20350.4 STA_VDBB.scala 260:29:@20589.4 STA_VDBB.scala 260:29:@20614.4 STA_VDBB.scala 260:29:@20853.4 STA_VDBB.scala 260:29:@20878.4 STA_VDBB.scala 260:29:@21117.4 STA_VDBB.scala 260:29:@21142.4 STA_VDBB.scala 339:29:@22101.4 STA_VDBB.scala 339:29:@22126.4 STA_VDBB.scala 339:29:@22893.4 STA_VDBB.scala 339:29:@22918.4 STA_VDBB.scala 339:29:@23685.4 STA_VDBB.scala 339:29:@23710.4 STA_VDBB.scala 339:29:@24477.4 STA_VDBB.scala 339:29:@24502.4 STA_VDBB.scala 339:29:@25269.4 STA_VDBB.scala 339:29:@25294.4 STA_VDBB.scala 339:29:@26061.4 STA_VDBB.scala 339:29:@26086.4 STA_VDBB.scala 339:29:@26853.4 STA_VDBB.scala 339:29:@26878.4 STA_VDBB.scala 339:29:@27645.4 STA_VDBB.scala 339:29:@27670.4]
  assign ffb1_io_in_tag_2_5 = S8DP1_14_io_out_tag_5; // @[STA_VDBB.scala 108:23:@10233.4 STA_VDBB.scala 127:29:@10438.4 STA_VDBB.scala 127:29:@10463.4 STA_VDBB.scala 127:29:@10702.4 STA_VDBB.scala 127:29:@10727.4 STA_VDBB.scala 127:29:@10966.4 STA_VDBB.scala 127:29:@10991.4 STA_VDBB.scala 127:29:@11230.4 STA_VDBB.scala 127:29:@11255.4 STA_VDBB.scala 127:29:@11494.4 STA_VDBB.scala 127:29:@11519.4 STA_VDBB.scala 127:29:@11758.4 STA_VDBB.scala 127:29:@11783.4 STA_VDBB.scala 127:29:@12022.4 STA_VDBB.scala 127:29:@12047.4 STA_VDBB.scala 127:29:@12286.4 STA_VDBB.scala 127:29:@12311.4 STA_VDBB.scala 207:29:@13270.4 STA_VDBB.scala 207:29:@13295.4 STA_VDBB.scala 207:29:@14062.4 STA_VDBB.scala 207:29:@14087.4 STA_VDBB.scala 207:29:@14854.4 STA_VDBB.scala 207:29:@14879.4 STA_VDBB.scala 207:29:@15646.4 STA_VDBB.scala 207:29:@15671.4 STA_VDBB.scala 207:29:@16438.4 STA_VDBB.scala 207:29:@16463.4 STA_VDBB.scala 207:29:@17230.4 STA_VDBB.scala 207:29:@17255.4 STA_VDBB.scala 207:29:@18022.4 STA_VDBB.scala 207:29:@18047.4 STA_VDBB.scala 207:29:@18814.4 STA_VDBB.scala 207:29:@18839.4 STA_VDBB.scala 241:23:@19065.4 STA_VDBB.scala 260:29:@19270.4 STA_VDBB.scala 260:29:@19295.4 STA_VDBB.scala 260:29:@19534.4 STA_VDBB.scala 260:29:@19559.4 STA_VDBB.scala 260:29:@19798.4 STA_VDBB.scala 260:29:@19823.4 STA_VDBB.scala 260:29:@20062.4 STA_VDBB.scala 260:29:@20087.4 STA_VDBB.scala 260:29:@20326.4 STA_VDBB.scala 260:29:@20351.4 STA_VDBB.scala 260:29:@20590.4 STA_VDBB.scala 260:29:@20615.4 STA_VDBB.scala 260:29:@20854.4 STA_VDBB.scala 260:29:@20879.4 STA_VDBB.scala 260:29:@21118.4 STA_VDBB.scala 260:29:@21143.4 STA_VDBB.scala 339:29:@22102.4 STA_VDBB.scala 339:29:@22127.4 STA_VDBB.scala 339:29:@22894.4 STA_VDBB.scala 339:29:@22919.4 STA_VDBB.scala 339:29:@23686.4 STA_VDBB.scala 339:29:@23711.4 STA_VDBB.scala 339:29:@24478.4 STA_VDBB.scala 339:29:@24503.4 STA_VDBB.scala 339:29:@25270.4 STA_VDBB.scala 339:29:@25295.4 STA_VDBB.scala 339:29:@26062.4 STA_VDBB.scala 339:29:@26087.4 STA_VDBB.scala 339:29:@26854.4 STA_VDBB.scala 339:29:@26879.4 STA_VDBB.scala 339:29:@27646.4 STA_VDBB.scala 339:29:@27671.4]
  assign ffb1_io_in_tag_2_6 = S8DP1_14_io_out_tag_6; // @[STA_VDBB.scala 108:23:@10234.4 STA_VDBB.scala 127:29:@10439.4 STA_VDBB.scala 127:29:@10464.4 STA_VDBB.scala 127:29:@10703.4 STA_VDBB.scala 127:29:@10728.4 STA_VDBB.scala 127:29:@10967.4 STA_VDBB.scala 127:29:@10992.4 STA_VDBB.scala 127:29:@11231.4 STA_VDBB.scala 127:29:@11256.4 STA_VDBB.scala 127:29:@11495.4 STA_VDBB.scala 127:29:@11520.4 STA_VDBB.scala 127:29:@11759.4 STA_VDBB.scala 127:29:@11784.4 STA_VDBB.scala 127:29:@12023.4 STA_VDBB.scala 127:29:@12048.4 STA_VDBB.scala 127:29:@12287.4 STA_VDBB.scala 127:29:@12312.4 STA_VDBB.scala 207:29:@13271.4 STA_VDBB.scala 207:29:@13296.4 STA_VDBB.scala 207:29:@14063.4 STA_VDBB.scala 207:29:@14088.4 STA_VDBB.scala 207:29:@14855.4 STA_VDBB.scala 207:29:@14880.4 STA_VDBB.scala 207:29:@15647.4 STA_VDBB.scala 207:29:@15672.4 STA_VDBB.scala 207:29:@16439.4 STA_VDBB.scala 207:29:@16464.4 STA_VDBB.scala 207:29:@17231.4 STA_VDBB.scala 207:29:@17256.4 STA_VDBB.scala 207:29:@18023.4 STA_VDBB.scala 207:29:@18048.4 STA_VDBB.scala 207:29:@18815.4 STA_VDBB.scala 207:29:@18840.4 STA_VDBB.scala 241:23:@19066.4 STA_VDBB.scala 260:29:@19271.4 STA_VDBB.scala 260:29:@19296.4 STA_VDBB.scala 260:29:@19535.4 STA_VDBB.scala 260:29:@19560.4 STA_VDBB.scala 260:29:@19799.4 STA_VDBB.scala 260:29:@19824.4 STA_VDBB.scala 260:29:@20063.4 STA_VDBB.scala 260:29:@20088.4 STA_VDBB.scala 260:29:@20327.4 STA_VDBB.scala 260:29:@20352.4 STA_VDBB.scala 260:29:@20591.4 STA_VDBB.scala 260:29:@20616.4 STA_VDBB.scala 260:29:@20855.4 STA_VDBB.scala 260:29:@20880.4 STA_VDBB.scala 260:29:@21119.4 STA_VDBB.scala 260:29:@21144.4 STA_VDBB.scala 339:29:@22103.4 STA_VDBB.scala 339:29:@22128.4 STA_VDBB.scala 339:29:@22895.4 STA_VDBB.scala 339:29:@22920.4 STA_VDBB.scala 339:29:@23687.4 STA_VDBB.scala 339:29:@23712.4 STA_VDBB.scala 339:29:@24479.4 STA_VDBB.scala 339:29:@24504.4 STA_VDBB.scala 339:29:@25271.4 STA_VDBB.scala 339:29:@25296.4 STA_VDBB.scala 339:29:@26063.4 STA_VDBB.scala 339:29:@26088.4 STA_VDBB.scala 339:29:@26855.4 STA_VDBB.scala 339:29:@26880.4 STA_VDBB.scala 339:29:@27647.4 STA_VDBB.scala 339:29:@27672.4]
  assign ffb1_io_in_tag_2_7 = S8DP1_14_io_out_tag_7; // @[STA_VDBB.scala 108:23:@10235.4 STA_VDBB.scala 127:29:@10440.4 STA_VDBB.scala 127:29:@10465.4 STA_VDBB.scala 127:29:@10704.4 STA_VDBB.scala 127:29:@10729.4 STA_VDBB.scala 127:29:@10968.4 STA_VDBB.scala 127:29:@10993.4 STA_VDBB.scala 127:29:@11232.4 STA_VDBB.scala 127:29:@11257.4 STA_VDBB.scala 127:29:@11496.4 STA_VDBB.scala 127:29:@11521.4 STA_VDBB.scala 127:29:@11760.4 STA_VDBB.scala 127:29:@11785.4 STA_VDBB.scala 127:29:@12024.4 STA_VDBB.scala 127:29:@12049.4 STA_VDBB.scala 127:29:@12288.4 STA_VDBB.scala 127:29:@12313.4 STA_VDBB.scala 207:29:@13272.4 STA_VDBB.scala 207:29:@13297.4 STA_VDBB.scala 207:29:@14064.4 STA_VDBB.scala 207:29:@14089.4 STA_VDBB.scala 207:29:@14856.4 STA_VDBB.scala 207:29:@14881.4 STA_VDBB.scala 207:29:@15648.4 STA_VDBB.scala 207:29:@15673.4 STA_VDBB.scala 207:29:@16440.4 STA_VDBB.scala 207:29:@16465.4 STA_VDBB.scala 207:29:@17232.4 STA_VDBB.scala 207:29:@17257.4 STA_VDBB.scala 207:29:@18024.4 STA_VDBB.scala 207:29:@18049.4 STA_VDBB.scala 207:29:@18816.4 STA_VDBB.scala 207:29:@18841.4 STA_VDBB.scala 241:23:@19067.4 STA_VDBB.scala 260:29:@19272.4 STA_VDBB.scala 260:29:@19297.4 STA_VDBB.scala 260:29:@19536.4 STA_VDBB.scala 260:29:@19561.4 STA_VDBB.scala 260:29:@19800.4 STA_VDBB.scala 260:29:@19825.4 STA_VDBB.scala 260:29:@20064.4 STA_VDBB.scala 260:29:@20089.4 STA_VDBB.scala 260:29:@20328.4 STA_VDBB.scala 260:29:@20353.4 STA_VDBB.scala 260:29:@20592.4 STA_VDBB.scala 260:29:@20617.4 STA_VDBB.scala 260:29:@20856.4 STA_VDBB.scala 260:29:@20881.4 STA_VDBB.scala 260:29:@21120.4 STA_VDBB.scala 260:29:@21145.4 STA_VDBB.scala 339:29:@22104.4 STA_VDBB.scala 339:29:@22129.4 STA_VDBB.scala 339:29:@22896.4 STA_VDBB.scala 339:29:@22921.4 STA_VDBB.scala 339:29:@23688.4 STA_VDBB.scala 339:29:@23713.4 STA_VDBB.scala 339:29:@24480.4 STA_VDBB.scala 339:29:@24505.4 STA_VDBB.scala 339:29:@25272.4 STA_VDBB.scala 339:29:@25297.4 STA_VDBB.scala 339:29:@26064.4 STA_VDBB.scala 339:29:@26089.4 STA_VDBB.scala 339:29:@26856.4 STA_VDBB.scala 339:29:@26881.4 STA_VDBB.scala 339:29:@27648.4 STA_VDBB.scala 339:29:@27673.4]
  assign ffb1_io_in_tag_3_0 = S8DP1_15_io_out_tag_0; // @[STA_VDBB.scala 108:23:@10252.4 STA_VDBB.scala 127:29:@10499.4 STA_VDBB.scala 127:29:@10524.4 STA_VDBB.scala 127:29:@10763.4 STA_VDBB.scala 127:29:@10788.4 STA_VDBB.scala 127:29:@11027.4 STA_VDBB.scala 127:29:@11052.4 STA_VDBB.scala 127:29:@11291.4 STA_VDBB.scala 127:29:@11316.4 STA_VDBB.scala 127:29:@11555.4 STA_VDBB.scala 127:29:@11580.4 STA_VDBB.scala 127:29:@11819.4 STA_VDBB.scala 127:29:@11844.4 STA_VDBB.scala 127:29:@12083.4 STA_VDBB.scala 127:29:@12108.4 STA_VDBB.scala 127:29:@12347.4 STA_VDBB.scala 127:29:@12372.4 STA_VDBB.scala 207:29:@13331.4 STA_VDBB.scala 207:29:@13356.4 STA_VDBB.scala 207:29:@14123.4 STA_VDBB.scala 207:29:@14148.4 STA_VDBB.scala 207:29:@14915.4 STA_VDBB.scala 207:29:@14940.4 STA_VDBB.scala 207:29:@15707.4 STA_VDBB.scala 207:29:@15732.4 STA_VDBB.scala 207:29:@16499.4 STA_VDBB.scala 207:29:@16524.4 STA_VDBB.scala 207:29:@17291.4 STA_VDBB.scala 207:29:@17316.4 STA_VDBB.scala 207:29:@18083.4 STA_VDBB.scala 207:29:@18108.4 STA_VDBB.scala 207:29:@18875.4 STA_VDBB.scala 207:29:@18900.4 STA_VDBB.scala 241:23:@19084.4 STA_VDBB.scala 260:29:@19331.4 STA_VDBB.scala 260:29:@19356.4 STA_VDBB.scala 260:29:@19595.4 STA_VDBB.scala 260:29:@19620.4 STA_VDBB.scala 260:29:@19859.4 STA_VDBB.scala 260:29:@19884.4 STA_VDBB.scala 260:29:@20123.4 STA_VDBB.scala 260:29:@20148.4 STA_VDBB.scala 260:29:@20387.4 STA_VDBB.scala 260:29:@20412.4 STA_VDBB.scala 260:29:@20651.4 STA_VDBB.scala 260:29:@20676.4 STA_VDBB.scala 260:29:@20915.4 STA_VDBB.scala 260:29:@20940.4 STA_VDBB.scala 260:29:@21179.4 STA_VDBB.scala 260:29:@21204.4 STA_VDBB.scala 339:29:@22163.4 STA_VDBB.scala 339:29:@22188.4 STA_VDBB.scala 339:29:@22955.4 STA_VDBB.scala 339:29:@22980.4 STA_VDBB.scala 339:29:@23747.4 STA_VDBB.scala 339:29:@23772.4 STA_VDBB.scala 339:29:@24539.4 STA_VDBB.scala 339:29:@24564.4 STA_VDBB.scala 339:29:@25331.4 STA_VDBB.scala 339:29:@25356.4 STA_VDBB.scala 339:29:@26123.4 STA_VDBB.scala 339:29:@26148.4 STA_VDBB.scala 339:29:@26915.4 STA_VDBB.scala 339:29:@26940.4 STA_VDBB.scala 339:29:@27707.4 STA_VDBB.scala 339:29:@27732.4]
  assign ffb1_io_in_tag_3_1 = S8DP1_15_io_out_tag_1; // @[STA_VDBB.scala 108:23:@10253.4 STA_VDBB.scala 127:29:@10500.4 STA_VDBB.scala 127:29:@10525.4 STA_VDBB.scala 127:29:@10764.4 STA_VDBB.scala 127:29:@10789.4 STA_VDBB.scala 127:29:@11028.4 STA_VDBB.scala 127:29:@11053.4 STA_VDBB.scala 127:29:@11292.4 STA_VDBB.scala 127:29:@11317.4 STA_VDBB.scala 127:29:@11556.4 STA_VDBB.scala 127:29:@11581.4 STA_VDBB.scala 127:29:@11820.4 STA_VDBB.scala 127:29:@11845.4 STA_VDBB.scala 127:29:@12084.4 STA_VDBB.scala 127:29:@12109.4 STA_VDBB.scala 127:29:@12348.4 STA_VDBB.scala 127:29:@12373.4 STA_VDBB.scala 207:29:@13332.4 STA_VDBB.scala 207:29:@13357.4 STA_VDBB.scala 207:29:@14124.4 STA_VDBB.scala 207:29:@14149.4 STA_VDBB.scala 207:29:@14916.4 STA_VDBB.scala 207:29:@14941.4 STA_VDBB.scala 207:29:@15708.4 STA_VDBB.scala 207:29:@15733.4 STA_VDBB.scala 207:29:@16500.4 STA_VDBB.scala 207:29:@16525.4 STA_VDBB.scala 207:29:@17292.4 STA_VDBB.scala 207:29:@17317.4 STA_VDBB.scala 207:29:@18084.4 STA_VDBB.scala 207:29:@18109.4 STA_VDBB.scala 207:29:@18876.4 STA_VDBB.scala 207:29:@18901.4 STA_VDBB.scala 241:23:@19085.4 STA_VDBB.scala 260:29:@19332.4 STA_VDBB.scala 260:29:@19357.4 STA_VDBB.scala 260:29:@19596.4 STA_VDBB.scala 260:29:@19621.4 STA_VDBB.scala 260:29:@19860.4 STA_VDBB.scala 260:29:@19885.4 STA_VDBB.scala 260:29:@20124.4 STA_VDBB.scala 260:29:@20149.4 STA_VDBB.scala 260:29:@20388.4 STA_VDBB.scala 260:29:@20413.4 STA_VDBB.scala 260:29:@20652.4 STA_VDBB.scala 260:29:@20677.4 STA_VDBB.scala 260:29:@20916.4 STA_VDBB.scala 260:29:@20941.4 STA_VDBB.scala 260:29:@21180.4 STA_VDBB.scala 260:29:@21205.4 STA_VDBB.scala 339:29:@22164.4 STA_VDBB.scala 339:29:@22189.4 STA_VDBB.scala 339:29:@22956.4 STA_VDBB.scala 339:29:@22981.4 STA_VDBB.scala 339:29:@23748.4 STA_VDBB.scala 339:29:@23773.4 STA_VDBB.scala 339:29:@24540.4 STA_VDBB.scala 339:29:@24565.4 STA_VDBB.scala 339:29:@25332.4 STA_VDBB.scala 339:29:@25357.4 STA_VDBB.scala 339:29:@26124.4 STA_VDBB.scala 339:29:@26149.4 STA_VDBB.scala 339:29:@26916.4 STA_VDBB.scala 339:29:@26941.4 STA_VDBB.scala 339:29:@27708.4 STA_VDBB.scala 339:29:@27733.4]
  assign ffb1_io_in_tag_3_2 = S8DP1_15_io_out_tag_2; // @[STA_VDBB.scala 108:23:@10254.4 STA_VDBB.scala 127:29:@10501.4 STA_VDBB.scala 127:29:@10526.4 STA_VDBB.scala 127:29:@10765.4 STA_VDBB.scala 127:29:@10790.4 STA_VDBB.scala 127:29:@11029.4 STA_VDBB.scala 127:29:@11054.4 STA_VDBB.scala 127:29:@11293.4 STA_VDBB.scala 127:29:@11318.4 STA_VDBB.scala 127:29:@11557.4 STA_VDBB.scala 127:29:@11582.4 STA_VDBB.scala 127:29:@11821.4 STA_VDBB.scala 127:29:@11846.4 STA_VDBB.scala 127:29:@12085.4 STA_VDBB.scala 127:29:@12110.4 STA_VDBB.scala 127:29:@12349.4 STA_VDBB.scala 127:29:@12374.4 STA_VDBB.scala 207:29:@13333.4 STA_VDBB.scala 207:29:@13358.4 STA_VDBB.scala 207:29:@14125.4 STA_VDBB.scala 207:29:@14150.4 STA_VDBB.scala 207:29:@14917.4 STA_VDBB.scala 207:29:@14942.4 STA_VDBB.scala 207:29:@15709.4 STA_VDBB.scala 207:29:@15734.4 STA_VDBB.scala 207:29:@16501.4 STA_VDBB.scala 207:29:@16526.4 STA_VDBB.scala 207:29:@17293.4 STA_VDBB.scala 207:29:@17318.4 STA_VDBB.scala 207:29:@18085.4 STA_VDBB.scala 207:29:@18110.4 STA_VDBB.scala 207:29:@18877.4 STA_VDBB.scala 207:29:@18902.4 STA_VDBB.scala 241:23:@19086.4 STA_VDBB.scala 260:29:@19333.4 STA_VDBB.scala 260:29:@19358.4 STA_VDBB.scala 260:29:@19597.4 STA_VDBB.scala 260:29:@19622.4 STA_VDBB.scala 260:29:@19861.4 STA_VDBB.scala 260:29:@19886.4 STA_VDBB.scala 260:29:@20125.4 STA_VDBB.scala 260:29:@20150.4 STA_VDBB.scala 260:29:@20389.4 STA_VDBB.scala 260:29:@20414.4 STA_VDBB.scala 260:29:@20653.4 STA_VDBB.scala 260:29:@20678.4 STA_VDBB.scala 260:29:@20917.4 STA_VDBB.scala 260:29:@20942.4 STA_VDBB.scala 260:29:@21181.4 STA_VDBB.scala 260:29:@21206.4 STA_VDBB.scala 339:29:@22165.4 STA_VDBB.scala 339:29:@22190.4 STA_VDBB.scala 339:29:@22957.4 STA_VDBB.scala 339:29:@22982.4 STA_VDBB.scala 339:29:@23749.4 STA_VDBB.scala 339:29:@23774.4 STA_VDBB.scala 339:29:@24541.4 STA_VDBB.scala 339:29:@24566.4 STA_VDBB.scala 339:29:@25333.4 STA_VDBB.scala 339:29:@25358.4 STA_VDBB.scala 339:29:@26125.4 STA_VDBB.scala 339:29:@26150.4 STA_VDBB.scala 339:29:@26917.4 STA_VDBB.scala 339:29:@26942.4 STA_VDBB.scala 339:29:@27709.4 STA_VDBB.scala 339:29:@27734.4]
  assign ffb1_io_in_tag_3_3 = S8DP1_15_io_out_tag_3; // @[STA_VDBB.scala 108:23:@10255.4 STA_VDBB.scala 127:29:@10502.4 STA_VDBB.scala 127:29:@10527.4 STA_VDBB.scala 127:29:@10766.4 STA_VDBB.scala 127:29:@10791.4 STA_VDBB.scala 127:29:@11030.4 STA_VDBB.scala 127:29:@11055.4 STA_VDBB.scala 127:29:@11294.4 STA_VDBB.scala 127:29:@11319.4 STA_VDBB.scala 127:29:@11558.4 STA_VDBB.scala 127:29:@11583.4 STA_VDBB.scala 127:29:@11822.4 STA_VDBB.scala 127:29:@11847.4 STA_VDBB.scala 127:29:@12086.4 STA_VDBB.scala 127:29:@12111.4 STA_VDBB.scala 127:29:@12350.4 STA_VDBB.scala 127:29:@12375.4 STA_VDBB.scala 207:29:@13334.4 STA_VDBB.scala 207:29:@13359.4 STA_VDBB.scala 207:29:@14126.4 STA_VDBB.scala 207:29:@14151.4 STA_VDBB.scala 207:29:@14918.4 STA_VDBB.scala 207:29:@14943.4 STA_VDBB.scala 207:29:@15710.4 STA_VDBB.scala 207:29:@15735.4 STA_VDBB.scala 207:29:@16502.4 STA_VDBB.scala 207:29:@16527.4 STA_VDBB.scala 207:29:@17294.4 STA_VDBB.scala 207:29:@17319.4 STA_VDBB.scala 207:29:@18086.4 STA_VDBB.scala 207:29:@18111.4 STA_VDBB.scala 207:29:@18878.4 STA_VDBB.scala 207:29:@18903.4 STA_VDBB.scala 241:23:@19087.4 STA_VDBB.scala 260:29:@19334.4 STA_VDBB.scala 260:29:@19359.4 STA_VDBB.scala 260:29:@19598.4 STA_VDBB.scala 260:29:@19623.4 STA_VDBB.scala 260:29:@19862.4 STA_VDBB.scala 260:29:@19887.4 STA_VDBB.scala 260:29:@20126.4 STA_VDBB.scala 260:29:@20151.4 STA_VDBB.scala 260:29:@20390.4 STA_VDBB.scala 260:29:@20415.4 STA_VDBB.scala 260:29:@20654.4 STA_VDBB.scala 260:29:@20679.4 STA_VDBB.scala 260:29:@20918.4 STA_VDBB.scala 260:29:@20943.4 STA_VDBB.scala 260:29:@21182.4 STA_VDBB.scala 260:29:@21207.4 STA_VDBB.scala 339:29:@22166.4 STA_VDBB.scala 339:29:@22191.4 STA_VDBB.scala 339:29:@22958.4 STA_VDBB.scala 339:29:@22983.4 STA_VDBB.scala 339:29:@23750.4 STA_VDBB.scala 339:29:@23775.4 STA_VDBB.scala 339:29:@24542.4 STA_VDBB.scala 339:29:@24567.4 STA_VDBB.scala 339:29:@25334.4 STA_VDBB.scala 339:29:@25359.4 STA_VDBB.scala 339:29:@26126.4 STA_VDBB.scala 339:29:@26151.4 STA_VDBB.scala 339:29:@26918.4 STA_VDBB.scala 339:29:@26943.4 STA_VDBB.scala 339:29:@27710.4 STA_VDBB.scala 339:29:@27735.4]
  assign ffb1_io_in_tag_3_4 = S8DP1_15_io_out_tag_4; // @[STA_VDBB.scala 108:23:@10256.4 STA_VDBB.scala 127:29:@10503.4 STA_VDBB.scala 127:29:@10528.4 STA_VDBB.scala 127:29:@10767.4 STA_VDBB.scala 127:29:@10792.4 STA_VDBB.scala 127:29:@11031.4 STA_VDBB.scala 127:29:@11056.4 STA_VDBB.scala 127:29:@11295.4 STA_VDBB.scala 127:29:@11320.4 STA_VDBB.scala 127:29:@11559.4 STA_VDBB.scala 127:29:@11584.4 STA_VDBB.scala 127:29:@11823.4 STA_VDBB.scala 127:29:@11848.4 STA_VDBB.scala 127:29:@12087.4 STA_VDBB.scala 127:29:@12112.4 STA_VDBB.scala 127:29:@12351.4 STA_VDBB.scala 127:29:@12376.4 STA_VDBB.scala 207:29:@13335.4 STA_VDBB.scala 207:29:@13360.4 STA_VDBB.scala 207:29:@14127.4 STA_VDBB.scala 207:29:@14152.4 STA_VDBB.scala 207:29:@14919.4 STA_VDBB.scala 207:29:@14944.4 STA_VDBB.scala 207:29:@15711.4 STA_VDBB.scala 207:29:@15736.4 STA_VDBB.scala 207:29:@16503.4 STA_VDBB.scala 207:29:@16528.4 STA_VDBB.scala 207:29:@17295.4 STA_VDBB.scala 207:29:@17320.4 STA_VDBB.scala 207:29:@18087.4 STA_VDBB.scala 207:29:@18112.4 STA_VDBB.scala 207:29:@18879.4 STA_VDBB.scala 207:29:@18904.4 STA_VDBB.scala 241:23:@19088.4 STA_VDBB.scala 260:29:@19335.4 STA_VDBB.scala 260:29:@19360.4 STA_VDBB.scala 260:29:@19599.4 STA_VDBB.scala 260:29:@19624.4 STA_VDBB.scala 260:29:@19863.4 STA_VDBB.scala 260:29:@19888.4 STA_VDBB.scala 260:29:@20127.4 STA_VDBB.scala 260:29:@20152.4 STA_VDBB.scala 260:29:@20391.4 STA_VDBB.scala 260:29:@20416.4 STA_VDBB.scala 260:29:@20655.4 STA_VDBB.scala 260:29:@20680.4 STA_VDBB.scala 260:29:@20919.4 STA_VDBB.scala 260:29:@20944.4 STA_VDBB.scala 260:29:@21183.4 STA_VDBB.scala 260:29:@21208.4 STA_VDBB.scala 339:29:@22167.4 STA_VDBB.scala 339:29:@22192.4 STA_VDBB.scala 339:29:@22959.4 STA_VDBB.scala 339:29:@22984.4 STA_VDBB.scala 339:29:@23751.4 STA_VDBB.scala 339:29:@23776.4 STA_VDBB.scala 339:29:@24543.4 STA_VDBB.scala 339:29:@24568.4 STA_VDBB.scala 339:29:@25335.4 STA_VDBB.scala 339:29:@25360.4 STA_VDBB.scala 339:29:@26127.4 STA_VDBB.scala 339:29:@26152.4 STA_VDBB.scala 339:29:@26919.4 STA_VDBB.scala 339:29:@26944.4 STA_VDBB.scala 339:29:@27711.4 STA_VDBB.scala 339:29:@27736.4]
  assign ffb1_io_in_tag_3_5 = S8DP1_15_io_out_tag_5; // @[STA_VDBB.scala 108:23:@10257.4 STA_VDBB.scala 127:29:@10504.4 STA_VDBB.scala 127:29:@10529.4 STA_VDBB.scala 127:29:@10768.4 STA_VDBB.scala 127:29:@10793.4 STA_VDBB.scala 127:29:@11032.4 STA_VDBB.scala 127:29:@11057.4 STA_VDBB.scala 127:29:@11296.4 STA_VDBB.scala 127:29:@11321.4 STA_VDBB.scala 127:29:@11560.4 STA_VDBB.scala 127:29:@11585.4 STA_VDBB.scala 127:29:@11824.4 STA_VDBB.scala 127:29:@11849.4 STA_VDBB.scala 127:29:@12088.4 STA_VDBB.scala 127:29:@12113.4 STA_VDBB.scala 127:29:@12352.4 STA_VDBB.scala 127:29:@12377.4 STA_VDBB.scala 207:29:@13336.4 STA_VDBB.scala 207:29:@13361.4 STA_VDBB.scala 207:29:@14128.4 STA_VDBB.scala 207:29:@14153.4 STA_VDBB.scala 207:29:@14920.4 STA_VDBB.scala 207:29:@14945.4 STA_VDBB.scala 207:29:@15712.4 STA_VDBB.scala 207:29:@15737.4 STA_VDBB.scala 207:29:@16504.4 STA_VDBB.scala 207:29:@16529.4 STA_VDBB.scala 207:29:@17296.4 STA_VDBB.scala 207:29:@17321.4 STA_VDBB.scala 207:29:@18088.4 STA_VDBB.scala 207:29:@18113.4 STA_VDBB.scala 207:29:@18880.4 STA_VDBB.scala 207:29:@18905.4 STA_VDBB.scala 241:23:@19089.4 STA_VDBB.scala 260:29:@19336.4 STA_VDBB.scala 260:29:@19361.4 STA_VDBB.scala 260:29:@19600.4 STA_VDBB.scala 260:29:@19625.4 STA_VDBB.scala 260:29:@19864.4 STA_VDBB.scala 260:29:@19889.4 STA_VDBB.scala 260:29:@20128.4 STA_VDBB.scala 260:29:@20153.4 STA_VDBB.scala 260:29:@20392.4 STA_VDBB.scala 260:29:@20417.4 STA_VDBB.scala 260:29:@20656.4 STA_VDBB.scala 260:29:@20681.4 STA_VDBB.scala 260:29:@20920.4 STA_VDBB.scala 260:29:@20945.4 STA_VDBB.scala 260:29:@21184.4 STA_VDBB.scala 260:29:@21209.4 STA_VDBB.scala 339:29:@22168.4 STA_VDBB.scala 339:29:@22193.4 STA_VDBB.scala 339:29:@22960.4 STA_VDBB.scala 339:29:@22985.4 STA_VDBB.scala 339:29:@23752.4 STA_VDBB.scala 339:29:@23777.4 STA_VDBB.scala 339:29:@24544.4 STA_VDBB.scala 339:29:@24569.4 STA_VDBB.scala 339:29:@25336.4 STA_VDBB.scala 339:29:@25361.4 STA_VDBB.scala 339:29:@26128.4 STA_VDBB.scala 339:29:@26153.4 STA_VDBB.scala 339:29:@26920.4 STA_VDBB.scala 339:29:@26945.4 STA_VDBB.scala 339:29:@27712.4 STA_VDBB.scala 339:29:@27737.4]
  assign ffb1_io_in_tag_3_6 = S8DP1_15_io_out_tag_6; // @[STA_VDBB.scala 108:23:@10258.4 STA_VDBB.scala 127:29:@10505.4 STA_VDBB.scala 127:29:@10530.4 STA_VDBB.scala 127:29:@10769.4 STA_VDBB.scala 127:29:@10794.4 STA_VDBB.scala 127:29:@11033.4 STA_VDBB.scala 127:29:@11058.4 STA_VDBB.scala 127:29:@11297.4 STA_VDBB.scala 127:29:@11322.4 STA_VDBB.scala 127:29:@11561.4 STA_VDBB.scala 127:29:@11586.4 STA_VDBB.scala 127:29:@11825.4 STA_VDBB.scala 127:29:@11850.4 STA_VDBB.scala 127:29:@12089.4 STA_VDBB.scala 127:29:@12114.4 STA_VDBB.scala 127:29:@12353.4 STA_VDBB.scala 127:29:@12378.4 STA_VDBB.scala 207:29:@13337.4 STA_VDBB.scala 207:29:@13362.4 STA_VDBB.scala 207:29:@14129.4 STA_VDBB.scala 207:29:@14154.4 STA_VDBB.scala 207:29:@14921.4 STA_VDBB.scala 207:29:@14946.4 STA_VDBB.scala 207:29:@15713.4 STA_VDBB.scala 207:29:@15738.4 STA_VDBB.scala 207:29:@16505.4 STA_VDBB.scala 207:29:@16530.4 STA_VDBB.scala 207:29:@17297.4 STA_VDBB.scala 207:29:@17322.4 STA_VDBB.scala 207:29:@18089.4 STA_VDBB.scala 207:29:@18114.4 STA_VDBB.scala 207:29:@18881.4 STA_VDBB.scala 207:29:@18906.4 STA_VDBB.scala 241:23:@19090.4 STA_VDBB.scala 260:29:@19337.4 STA_VDBB.scala 260:29:@19362.4 STA_VDBB.scala 260:29:@19601.4 STA_VDBB.scala 260:29:@19626.4 STA_VDBB.scala 260:29:@19865.4 STA_VDBB.scala 260:29:@19890.4 STA_VDBB.scala 260:29:@20129.4 STA_VDBB.scala 260:29:@20154.4 STA_VDBB.scala 260:29:@20393.4 STA_VDBB.scala 260:29:@20418.4 STA_VDBB.scala 260:29:@20657.4 STA_VDBB.scala 260:29:@20682.4 STA_VDBB.scala 260:29:@20921.4 STA_VDBB.scala 260:29:@20946.4 STA_VDBB.scala 260:29:@21185.4 STA_VDBB.scala 260:29:@21210.4 STA_VDBB.scala 339:29:@22169.4 STA_VDBB.scala 339:29:@22194.4 STA_VDBB.scala 339:29:@22961.4 STA_VDBB.scala 339:29:@22986.4 STA_VDBB.scala 339:29:@23753.4 STA_VDBB.scala 339:29:@23778.4 STA_VDBB.scala 339:29:@24545.4 STA_VDBB.scala 339:29:@24570.4 STA_VDBB.scala 339:29:@25337.4 STA_VDBB.scala 339:29:@25362.4 STA_VDBB.scala 339:29:@26129.4 STA_VDBB.scala 339:29:@26154.4 STA_VDBB.scala 339:29:@26921.4 STA_VDBB.scala 339:29:@26946.4 STA_VDBB.scala 339:29:@27713.4 STA_VDBB.scala 339:29:@27738.4]
  assign ffb1_io_in_tag_3_7 = S8DP1_15_io_out_tag_7; // @[STA_VDBB.scala 108:23:@10259.4 STA_VDBB.scala 127:29:@10506.4 STA_VDBB.scala 127:29:@10531.4 STA_VDBB.scala 127:29:@10770.4 STA_VDBB.scala 127:29:@10795.4 STA_VDBB.scala 127:29:@11034.4 STA_VDBB.scala 127:29:@11059.4 STA_VDBB.scala 127:29:@11298.4 STA_VDBB.scala 127:29:@11323.4 STA_VDBB.scala 127:29:@11562.4 STA_VDBB.scala 127:29:@11587.4 STA_VDBB.scala 127:29:@11826.4 STA_VDBB.scala 127:29:@11851.4 STA_VDBB.scala 127:29:@12090.4 STA_VDBB.scala 127:29:@12115.4 STA_VDBB.scala 127:29:@12354.4 STA_VDBB.scala 127:29:@12379.4 STA_VDBB.scala 207:29:@13338.4 STA_VDBB.scala 207:29:@13363.4 STA_VDBB.scala 207:29:@14130.4 STA_VDBB.scala 207:29:@14155.4 STA_VDBB.scala 207:29:@14922.4 STA_VDBB.scala 207:29:@14947.4 STA_VDBB.scala 207:29:@15714.4 STA_VDBB.scala 207:29:@15739.4 STA_VDBB.scala 207:29:@16506.4 STA_VDBB.scala 207:29:@16531.4 STA_VDBB.scala 207:29:@17298.4 STA_VDBB.scala 207:29:@17323.4 STA_VDBB.scala 207:29:@18090.4 STA_VDBB.scala 207:29:@18115.4 STA_VDBB.scala 207:29:@18882.4 STA_VDBB.scala 207:29:@18907.4 STA_VDBB.scala 241:23:@19091.4 STA_VDBB.scala 260:29:@19338.4 STA_VDBB.scala 260:29:@19363.4 STA_VDBB.scala 260:29:@19602.4 STA_VDBB.scala 260:29:@19627.4 STA_VDBB.scala 260:29:@19866.4 STA_VDBB.scala 260:29:@19891.4 STA_VDBB.scala 260:29:@20130.4 STA_VDBB.scala 260:29:@20155.4 STA_VDBB.scala 260:29:@20394.4 STA_VDBB.scala 260:29:@20419.4 STA_VDBB.scala 260:29:@20658.4 STA_VDBB.scala 260:29:@20683.4 STA_VDBB.scala 260:29:@20922.4 STA_VDBB.scala 260:29:@20947.4 STA_VDBB.scala 260:29:@21186.4 STA_VDBB.scala 260:29:@21211.4 STA_VDBB.scala 339:29:@22170.4 STA_VDBB.scala 339:29:@22195.4 STA_VDBB.scala 339:29:@22962.4 STA_VDBB.scala 339:29:@22987.4 STA_VDBB.scala 339:29:@23754.4 STA_VDBB.scala 339:29:@23779.4 STA_VDBB.scala 339:29:@24546.4 STA_VDBB.scala 339:29:@24571.4 STA_VDBB.scala 339:29:@25338.4 STA_VDBB.scala 339:29:@25363.4 STA_VDBB.scala 339:29:@26130.4 STA_VDBB.scala 339:29:@26155.4 STA_VDBB.scala 339:29:@26922.4 STA_VDBB.scala 339:29:@26947.4 STA_VDBB.scala 339:29:@27714.4 STA_VDBB.scala 339:29:@27739.4]
  assign ffb2_clock = clock; // @[:@9790.4]
  assign ffb2_reset = reset; // @[:@9791.4]
  assign ffb2_io_in_data_0_0 = io_in_B_4_8; // @[STA_VDBB.scala 153:29:@12384.4 STA_VDBB.scala 285:29:@21216.4]
  assign ffb2_io_in_data_0_1 = io_in_B_4_9; // @[STA_VDBB.scala 153:29:@12396.4 STA_VDBB.scala 285:29:@21228.4]
  assign ffb2_io_in_data_0_2 = io_in_B_4_10; // @[STA_VDBB.scala 153:29:@12408.4 STA_VDBB.scala 285:29:@21240.4]
  assign ffb2_io_in_data_0_3 = io_in_B_4_11; // @[STA_VDBB.scala 153:29:@12420.4 STA_VDBB.scala 285:29:@21252.4]
  assign ffb2_io_in_data_0_4 = io_in_B_4_12; // @[STA_VDBB.scala 153:29:@12432.4 STA_VDBB.scala 285:29:@21264.4]
  assign ffb2_io_in_data_0_5 = io_in_B_4_13; // @[STA_VDBB.scala 153:29:@12444.4 STA_VDBB.scala 285:29:@21276.4]
  assign ffb2_io_in_data_0_6 = io_in_B_4_14; // @[STA_VDBB.scala 153:29:@12456.4 STA_VDBB.scala 285:29:@21288.4]
  assign ffb2_io_in_data_0_7 = io_in_B_4_15; // @[STA_VDBB.scala 153:29:@12468.4 STA_VDBB.scala 285:29:@21300.4]
  assign ffb2_io_in_data_1_0 = io_in_B_5_8; // @[STA_VDBB.scala 153:29:@12386.4 STA_VDBB.scala 285:29:@21218.4]
  assign ffb2_io_in_data_1_1 = io_in_B_5_9; // @[STA_VDBB.scala 153:29:@12398.4 STA_VDBB.scala 285:29:@21230.4]
  assign ffb2_io_in_data_1_2 = io_in_B_5_10; // @[STA_VDBB.scala 153:29:@12410.4 STA_VDBB.scala 285:29:@21242.4]
  assign ffb2_io_in_data_1_3 = io_in_B_5_11; // @[STA_VDBB.scala 153:29:@12422.4 STA_VDBB.scala 285:29:@21254.4]
  assign ffb2_io_in_data_1_4 = io_in_B_5_12; // @[STA_VDBB.scala 153:29:@12434.4 STA_VDBB.scala 285:29:@21266.4]
  assign ffb2_io_in_data_1_5 = io_in_B_5_13; // @[STA_VDBB.scala 153:29:@12446.4 STA_VDBB.scala 285:29:@21278.4]
  assign ffb2_io_in_data_1_6 = io_in_B_5_14; // @[STA_VDBB.scala 153:29:@12458.4 STA_VDBB.scala 285:29:@21290.4]
  assign ffb2_io_in_data_1_7 = io_in_B_5_15; // @[STA_VDBB.scala 153:29:@12470.4 STA_VDBB.scala 285:29:@21302.4]
  assign ffb2_io_in_data_2_0 = io_in_B_6_8; // @[STA_VDBB.scala 153:29:@12388.4 STA_VDBB.scala 285:29:@21220.4]
  assign ffb2_io_in_data_2_1 = io_in_B_6_9; // @[STA_VDBB.scala 153:29:@12400.4 STA_VDBB.scala 285:29:@21232.4]
  assign ffb2_io_in_data_2_2 = io_in_B_6_10; // @[STA_VDBB.scala 153:29:@12412.4 STA_VDBB.scala 285:29:@21244.4]
  assign ffb2_io_in_data_2_3 = io_in_B_6_11; // @[STA_VDBB.scala 153:29:@12424.4 STA_VDBB.scala 285:29:@21256.4]
  assign ffb2_io_in_data_2_4 = io_in_B_6_12; // @[STA_VDBB.scala 153:29:@12436.4 STA_VDBB.scala 285:29:@21268.4]
  assign ffb2_io_in_data_2_5 = io_in_B_6_13; // @[STA_VDBB.scala 153:29:@12448.4 STA_VDBB.scala 285:29:@21280.4]
  assign ffb2_io_in_data_2_6 = io_in_B_6_14; // @[STA_VDBB.scala 153:29:@12460.4 STA_VDBB.scala 285:29:@21292.4]
  assign ffb2_io_in_data_2_7 = io_in_B_6_15; // @[STA_VDBB.scala 153:29:@12472.4 STA_VDBB.scala 285:29:@21304.4]
  assign ffb2_io_in_data_3_0 = io_in_B_7_8; // @[STA_VDBB.scala 153:29:@12390.4 STA_VDBB.scala 285:29:@21222.4]
  assign ffb2_io_in_data_3_1 = io_in_B_7_9; // @[STA_VDBB.scala 153:29:@12402.4 STA_VDBB.scala 285:29:@21234.4]
  assign ffb2_io_in_data_3_2 = io_in_B_7_10; // @[STA_VDBB.scala 153:29:@12414.4 STA_VDBB.scala 285:29:@21246.4]
  assign ffb2_io_in_data_3_3 = io_in_B_7_11; // @[STA_VDBB.scala 153:29:@12426.4 STA_VDBB.scala 285:29:@21258.4]
  assign ffb2_io_in_data_3_4 = io_in_B_7_12; // @[STA_VDBB.scala 153:29:@12438.4 STA_VDBB.scala 285:29:@21270.4]
  assign ffb2_io_in_data_3_5 = io_in_B_7_13; // @[STA_VDBB.scala 153:29:@12450.4 STA_VDBB.scala 285:29:@21282.4]
  assign ffb2_io_in_data_3_6 = io_in_B_7_14; // @[STA_VDBB.scala 153:29:@12462.4 STA_VDBB.scala 285:29:@21294.4]
  assign ffb2_io_in_data_3_7 = io_in_B_7_15; // @[STA_VDBB.scala 153:29:@12474.4 STA_VDBB.scala 285:29:@21306.4]
  assign ffb2_io_in_tag_0_0 = S8DP1_12_io_out_tag_0; // @[STA_VDBB.scala 161:23:@12484.4 STA_VDBB.scala 181:29:@12605.4 STA_VDBB.scala 181:29:@12630.4 STA_VDBB.scala 181:29:@13397.4 STA_VDBB.scala 181:29:@13422.4 STA_VDBB.scala 181:29:@14189.4 STA_VDBB.scala 181:29:@14214.4 STA_VDBB.scala 181:29:@14981.4 STA_VDBB.scala 181:29:@15006.4 STA_VDBB.scala 181:29:@15773.4 STA_VDBB.scala 181:29:@15798.4 STA_VDBB.scala 181:29:@16565.4 STA_VDBB.scala 181:29:@16590.4 STA_VDBB.scala 181:29:@17357.4 STA_VDBB.scala 181:29:@17382.4 STA_VDBB.scala 181:29:@18149.4 STA_VDBB.scala 181:29:@18174.4 STA_VDBB.scala 293:23:@21316.4 STA_VDBB.scala 313:29:@21437.4 STA_VDBB.scala 313:29:@21462.4 STA_VDBB.scala 313:29:@22229.4 STA_VDBB.scala 313:29:@22254.4 STA_VDBB.scala 313:29:@23021.4 STA_VDBB.scala 313:29:@23046.4 STA_VDBB.scala 313:29:@23813.4 STA_VDBB.scala 313:29:@23838.4 STA_VDBB.scala 313:29:@24605.4 STA_VDBB.scala 313:29:@24630.4 STA_VDBB.scala 313:29:@25397.4 STA_VDBB.scala 313:29:@25422.4 STA_VDBB.scala 313:29:@26189.4 STA_VDBB.scala 313:29:@26214.4 STA_VDBB.scala 313:29:@26981.4 STA_VDBB.scala 313:29:@27006.4]
  assign ffb2_io_in_tag_0_1 = S8DP1_12_io_out_tag_1; // @[STA_VDBB.scala 161:23:@12485.4 STA_VDBB.scala 181:29:@12606.4 STA_VDBB.scala 181:29:@12631.4 STA_VDBB.scala 181:29:@13398.4 STA_VDBB.scala 181:29:@13423.4 STA_VDBB.scala 181:29:@14190.4 STA_VDBB.scala 181:29:@14215.4 STA_VDBB.scala 181:29:@14982.4 STA_VDBB.scala 181:29:@15007.4 STA_VDBB.scala 181:29:@15774.4 STA_VDBB.scala 181:29:@15799.4 STA_VDBB.scala 181:29:@16566.4 STA_VDBB.scala 181:29:@16591.4 STA_VDBB.scala 181:29:@17358.4 STA_VDBB.scala 181:29:@17383.4 STA_VDBB.scala 181:29:@18150.4 STA_VDBB.scala 181:29:@18175.4 STA_VDBB.scala 293:23:@21317.4 STA_VDBB.scala 313:29:@21438.4 STA_VDBB.scala 313:29:@21463.4 STA_VDBB.scala 313:29:@22230.4 STA_VDBB.scala 313:29:@22255.4 STA_VDBB.scala 313:29:@23022.4 STA_VDBB.scala 313:29:@23047.4 STA_VDBB.scala 313:29:@23814.4 STA_VDBB.scala 313:29:@23839.4 STA_VDBB.scala 313:29:@24606.4 STA_VDBB.scala 313:29:@24631.4 STA_VDBB.scala 313:29:@25398.4 STA_VDBB.scala 313:29:@25423.4 STA_VDBB.scala 313:29:@26190.4 STA_VDBB.scala 313:29:@26215.4 STA_VDBB.scala 313:29:@26982.4 STA_VDBB.scala 313:29:@27007.4]
  assign ffb2_io_in_tag_0_2 = S8DP1_12_io_out_tag_2; // @[STA_VDBB.scala 161:23:@12486.4 STA_VDBB.scala 181:29:@12607.4 STA_VDBB.scala 181:29:@12632.4 STA_VDBB.scala 181:29:@13399.4 STA_VDBB.scala 181:29:@13424.4 STA_VDBB.scala 181:29:@14191.4 STA_VDBB.scala 181:29:@14216.4 STA_VDBB.scala 181:29:@14983.4 STA_VDBB.scala 181:29:@15008.4 STA_VDBB.scala 181:29:@15775.4 STA_VDBB.scala 181:29:@15800.4 STA_VDBB.scala 181:29:@16567.4 STA_VDBB.scala 181:29:@16592.4 STA_VDBB.scala 181:29:@17359.4 STA_VDBB.scala 181:29:@17384.4 STA_VDBB.scala 181:29:@18151.4 STA_VDBB.scala 181:29:@18176.4 STA_VDBB.scala 293:23:@21318.4 STA_VDBB.scala 313:29:@21439.4 STA_VDBB.scala 313:29:@21464.4 STA_VDBB.scala 313:29:@22231.4 STA_VDBB.scala 313:29:@22256.4 STA_VDBB.scala 313:29:@23023.4 STA_VDBB.scala 313:29:@23048.4 STA_VDBB.scala 313:29:@23815.4 STA_VDBB.scala 313:29:@23840.4 STA_VDBB.scala 313:29:@24607.4 STA_VDBB.scala 313:29:@24632.4 STA_VDBB.scala 313:29:@25399.4 STA_VDBB.scala 313:29:@25424.4 STA_VDBB.scala 313:29:@26191.4 STA_VDBB.scala 313:29:@26216.4 STA_VDBB.scala 313:29:@26983.4 STA_VDBB.scala 313:29:@27008.4]
  assign ffb2_io_in_tag_0_3 = S8DP1_12_io_out_tag_3; // @[STA_VDBB.scala 161:23:@12487.4 STA_VDBB.scala 181:29:@12608.4 STA_VDBB.scala 181:29:@12633.4 STA_VDBB.scala 181:29:@13400.4 STA_VDBB.scala 181:29:@13425.4 STA_VDBB.scala 181:29:@14192.4 STA_VDBB.scala 181:29:@14217.4 STA_VDBB.scala 181:29:@14984.4 STA_VDBB.scala 181:29:@15009.4 STA_VDBB.scala 181:29:@15776.4 STA_VDBB.scala 181:29:@15801.4 STA_VDBB.scala 181:29:@16568.4 STA_VDBB.scala 181:29:@16593.4 STA_VDBB.scala 181:29:@17360.4 STA_VDBB.scala 181:29:@17385.4 STA_VDBB.scala 181:29:@18152.4 STA_VDBB.scala 181:29:@18177.4 STA_VDBB.scala 293:23:@21319.4 STA_VDBB.scala 313:29:@21440.4 STA_VDBB.scala 313:29:@21465.4 STA_VDBB.scala 313:29:@22232.4 STA_VDBB.scala 313:29:@22257.4 STA_VDBB.scala 313:29:@23024.4 STA_VDBB.scala 313:29:@23049.4 STA_VDBB.scala 313:29:@23816.4 STA_VDBB.scala 313:29:@23841.4 STA_VDBB.scala 313:29:@24608.4 STA_VDBB.scala 313:29:@24633.4 STA_VDBB.scala 313:29:@25400.4 STA_VDBB.scala 313:29:@25425.4 STA_VDBB.scala 313:29:@26192.4 STA_VDBB.scala 313:29:@26217.4 STA_VDBB.scala 313:29:@26984.4 STA_VDBB.scala 313:29:@27009.4]
  assign ffb2_io_in_tag_0_4 = S8DP1_12_io_out_tag_4; // @[STA_VDBB.scala 161:23:@12488.4 STA_VDBB.scala 181:29:@12609.4 STA_VDBB.scala 181:29:@12634.4 STA_VDBB.scala 181:29:@13401.4 STA_VDBB.scala 181:29:@13426.4 STA_VDBB.scala 181:29:@14193.4 STA_VDBB.scala 181:29:@14218.4 STA_VDBB.scala 181:29:@14985.4 STA_VDBB.scala 181:29:@15010.4 STA_VDBB.scala 181:29:@15777.4 STA_VDBB.scala 181:29:@15802.4 STA_VDBB.scala 181:29:@16569.4 STA_VDBB.scala 181:29:@16594.4 STA_VDBB.scala 181:29:@17361.4 STA_VDBB.scala 181:29:@17386.4 STA_VDBB.scala 181:29:@18153.4 STA_VDBB.scala 181:29:@18178.4 STA_VDBB.scala 293:23:@21320.4 STA_VDBB.scala 313:29:@21441.4 STA_VDBB.scala 313:29:@21466.4 STA_VDBB.scala 313:29:@22233.4 STA_VDBB.scala 313:29:@22258.4 STA_VDBB.scala 313:29:@23025.4 STA_VDBB.scala 313:29:@23050.4 STA_VDBB.scala 313:29:@23817.4 STA_VDBB.scala 313:29:@23842.4 STA_VDBB.scala 313:29:@24609.4 STA_VDBB.scala 313:29:@24634.4 STA_VDBB.scala 313:29:@25401.4 STA_VDBB.scala 313:29:@25426.4 STA_VDBB.scala 313:29:@26193.4 STA_VDBB.scala 313:29:@26218.4 STA_VDBB.scala 313:29:@26985.4 STA_VDBB.scala 313:29:@27010.4]
  assign ffb2_io_in_tag_0_5 = S8DP1_12_io_out_tag_5; // @[STA_VDBB.scala 161:23:@12489.4 STA_VDBB.scala 181:29:@12610.4 STA_VDBB.scala 181:29:@12635.4 STA_VDBB.scala 181:29:@13402.4 STA_VDBB.scala 181:29:@13427.4 STA_VDBB.scala 181:29:@14194.4 STA_VDBB.scala 181:29:@14219.4 STA_VDBB.scala 181:29:@14986.4 STA_VDBB.scala 181:29:@15011.4 STA_VDBB.scala 181:29:@15778.4 STA_VDBB.scala 181:29:@15803.4 STA_VDBB.scala 181:29:@16570.4 STA_VDBB.scala 181:29:@16595.4 STA_VDBB.scala 181:29:@17362.4 STA_VDBB.scala 181:29:@17387.4 STA_VDBB.scala 181:29:@18154.4 STA_VDBB.scala 181:29:@18179.4 STA_VDBB.scala 293:23:@21321.4 STA_VDBB.scala 313:29:@21442.4 STA_VDBB.scala 313:29:@21467.4 STA_VDBB.scala 313:29:@22234.4 STA_VDBB.scala 313:29:@22259.4 STA_VDBB.scala 313:29:@23026.4 STA_VDBB.scala 313:29:@23051.4 STA_VDBB.scala 313:29:@23818.4 STA_VDBB.scala 313:29:@23843.4 STA_VDBB.scala 313:29:@24610.4 STA_VDBB.scala 313:29:@24635.4 STA_VDBB.scala 313:29:@25402.4 STA_VDBB.scala 313:29:@25427.4 STA_VDBB.scala 313:29:@26194.4 STA_VDBB.scala 313:29:@26219.4 STA_VDBB.scala 313:29:@26986.4 STA_VDBB.scala 313:29:@27011.4]
  assign ffb2_io_in_tag_0_6 = S8DP1_12_io_out_tag_6; // @[STA_VDBB.scala 161:23:@12490.4 STA_VDBB.scala 181:29:@12611.4 STA_VDBB.scala 181:29:@12636.4 STA_VDBB.scala 181:29:@13403.4 STA_VDBB.scala 181:29:@13428.4 STA_VDBB.scala 181:29:@14195.4 STA_VDBB.scala 181:29:@14220.4 STA_VDBB.scala 181:29:@14987.4 STA_VDBB.scala 181:29:@15012.4 STA_VDBB.scala 181:29:@15779.4 STA_VDBB.scala 181:29:@15804.4 STA_VDBB.scala 181:29:@16571.4 STA_VDBB.scala 181:29:@16596.4 STA_VDBB.scala 181:29:@17363.4 STA_VDBB.scala 181:29:@17388.4 STA_VDBB.scala 181:29:@18155.4 STA_VDBB.scala 181:29:@18180.4 STA_VDBB.scala 293:23:@21322.4 STA_VDBB.scala 313:29:@21443.4 STA_VDBB.scala 313:29:@21468.4 STA_VDBB.scala 313:29:@22235.4 STA_VDBB.scala 313:29:@22260.4 STA_VDBB.scala 313:29:@23027.4 STA_VDBB.scala 313:29:@23052.4 STA_VDBB.scala 313:29:@23819.4 STA_VDBB.scala 313:29:@23844.4 STA_VDBB.scala 313:29:@24611.4 STA_VDBB.scala 313:29:@24636.4 STA_VDBB.scala 313:29:@25403.4 STA_VDBB.scala 313:29:@25428.4 STA_VDBB.scala 313:29:@26195.4 STA_VDBB.scala 313:29:@26220.4 STA_VDBB.scala 313:29:@26987.4 STA_VDBB.scala 313:29:@27012.4]
  assign ffb2_io_in_tag_0_7 = S8DP1_12_io_out_tag_7; // @[STA_VDBB.scala 161:23:@12491.4 STA_VDBB.scala 181:29:@12612.4 STA_VDBB.scala 181:29:@12637.4 STA_VDBB.scala 181:29:@13404.4 STA_VDBB.scala 181:29:@13429.4 STA_VDBB.scala 181:29:@14196.4 STA_VDBB.scala 181:29:@14221.4 STA_VDBB.scala 181:29:@14988.4 STA_VDBB.scala 181:29:@15013.4 STA_VDBB.scala 181:29:@15780.4 STA_VDBB.scala 181:29:@15805.4 STA_VDBB.scala 181:29:@16572.4 STA_VDBB.scala 181:29:@16597.4 STA_VDBB.scala 181:29:@17364.4 STA_VDBB.scala 181:29:@17389.4 STA_VDBB.scala 181:29:@18156.4 STA_VDBB.scala 181:29:@18181.4 STA_VDBB.scala 293:23:@21323.4 STA_VDBB.scala 313:29:@21444.4 STA_VDBB.scala 313:29:@21469.4 STA_VDBB.scala 313:29:@22236.4 STA_VDBB.scala 313:29:@22261.4 STA_VDBB.scala 313:29:@23028.4 STA_VDBB.scala 313:29:@23053.4 STA_VDBB.scala 313:29:@23820.4 STA_VDBB.scala 313:29:@23845.4 STA_VDBB.scala 313:29:@24612.4 STA_VDBB.scala 313:29:@24637.4 STA_VDBB.scala 313:29:@25404.4 STA_VDBB.scala 313:29:@25429.4 STA_VDBB.scala 313:29:@26196.4 STA_VDBB.scala 313:29:@26221.4 STA_VDBB.scala 313:29:@26988.4 STA_VDBB.scala 313:29:@27013.4]
  assign ffb2_io_in_tag_1_0 = S8DP1_13_io_out_tag_0; // @[STA_VDBB.scala 161:23:@12508.4 STA_VDBB.scala 181:29:@12671.4 STA_VDBB.scala 181:29:@12696.4 STA_VDBB.scala 181:29:@13463.4 STA_VDBB.scala 181:29:@13488.4 STA_VDBB.scala 181:29:@14255.4 STA_VDBB.scala 181:29:@14280.4 STA_VDBB.scala 181:29:@15047.4 STA_VDBB.scala 181:29:@15072.4 STA_VDBB.scala 181:29:@15839.4 STA_VDBB.scala 181:29:@15864.4 STA_VDBB.scala 181:29:@16631.4 STA_VDBB.scala 181:29:@16656.4 STA_VDBB.scala 181:29:@17423.4 STA_VDBB.scala 181:29:@17448.4 STA_VDBB.scala 181:29:@18215.4 STA_VDBB.scala 181:29:@18240.4 STA_VDBB.scala 293:23:@21340.4 STA_VDBB.scala 313:29:@21503.4 STA_VDBB.scala 313:29:@21528.4 STA_VDBB.scala 313:29:@22295.4 STA_VDBB.scala 313:29:@22320.4 STA_VDBB.scala 313:29:@23087.4 STA_VDBB.scala 313:29:@23112.4 STA_VDBB.scala 313:29:@23879.4 STA_VDBB.scala 313:29:@23904.4 STA_VDBB.scala 313:29:@24671.4 STA_VDBB.scala 313:29:@24696.4 STA_VDBB.scala 313:29:@25463.4 STA_VDBB.scala 313:29:@25488.4 STA_VDBB.scala 313:29:@26255.4 STA_VDBB.scala 313:29:@26280.4 STA_VDBB.scala 313:29:@27047.4 STA_VDBB.scala 313:29:@27072.4]
  assign ffb2_io_in_tag_1_1 = S8DP1_13_io_out_tag_1; // @[STA_VDBB.scala 161:23:@12509.4 STA_VDBB.scala 181:29:@12672.4 STA_VDBB.scala 181:29:@12697.4 STA_VDBB.scala 181:29:@13464.4 STA_VDBB.scala 181:29:@13489.4 STA_VDBB.scala 181:29:@14256.4 STA_VDBB.scala 181:29:@14281.4 STA_VDBB.scala 181:29:@15048.4 STA_VDBB.scala 181:29:@15073.4 STA_VDBB.scala 181:29:@15840.4 STA_VDBB.scala 181:29:@15865.4 STA_VDBB.scala 181:29:@16632.4 STA_VDBB.scala 181:29:@16657.4 STA_VDBB.scala 181:29:@17424.4 STA_VDBB.scala 181:29:@17449.4 STA_VDBB.scala 181:29:@18216.4 STA_VDBB.scala 181:29:@18241.4 STA_VDBB.scala 293:23:@21341.4 STA_VDBB.scala 313:29:@21504.4 STA_VDBB.scala 313:29:@21529.4 STA_VDBB.scala 313:29:@22296.4 STA_VDBB.scala 313:29:@22321.4 STA_VDBB.scala 313:29:@23088.4 STA_VDBB.scala 313:29:@23113.4 STA_VDBB.scala 313:29:@23880.4 STA_VDBB.scala 313:29:@23905.4 STA_VDBB.scala 313:29:@24672.4 STA_VDBB.scala 313:29:@24697.4 STA_VDBB.scala 313:29:@25464.4 STA_VDBB.scala 313:29:@25489.4 STA_VDBB.scala 313:29:@26256.4 STA_VDBB.scala 313:29:@26281.4 STA_VDBB.scala 313:29:@27048.4 STA_VDBB.scala 313:29:@27073.4]
  assign ffb2_io_in_tag_1_2 = S8DP1_13_io_out_tag_2; // @[STA_VDBB.scala 161:23:@12510.4 STA_VDBB.scala 181:29:@12673.4 STA_VDBB.scala 181:29:@12698.4 STA_VDBB.scala 181:29:@13465.4 STA_VDBB.scala 181:29:@13490.4 STA_VDBB.scala 181:29:@14257.4 STA_VDBB.scala 181:29:@14282.4 STA_VDBB.scala 181:29:@15049.4 STA_VDBB.scala 181:29:@15074.4 STA_VDBB.scala 181:29:@15841.4 STA_VDBB.scala 181:29:@15866.4 STA_VDBB.scala 181:29:@16633.4 STA_VDBB.scala 181:29:@16658.4 STA_VDBB.scala 181:29:@17425.4 STA_VDBB.scala 181:29:@17450.4 STA_VDBB.scala 181:29:@18217.4 STA_VDBB.scala 181:29:@18242.4 STA_VDBB.scala 293:23:@21342.4 STA_VDBB.scala 313:29:@21505.4 STA_VDBB.scala 313:29:@21530.4 STA_VDBB.scala 313:29:@22297.4 STA_VDBB.scala 313:29:@22322.4 STA_VDBB.scala 313:29:@23089.4 STA_VDBB.scala 313:29:@23114.4 STA_VDBB.scala 313:29:@23881.4 STA_VDBB.scala 313:29:@23906.4 STA_VDBB.scala 313:29:@24673.4 STA_VDBB.scala 313:29:@24698.4 STA_VDBB.scala 313:29:@25465.4 STA_VDBB.scala 313:29:@25490.4 STA_VDBB.scala 313:29:@26257.4 STA_VDBB.scala 313:29:@26282.4 STA_VDBB.scala 313:29:@27049.4 STA_VDBB.scala 313:29:@27074.4]
  assign ffb2_io_in_tag_1_3 = S8DP1_13_io_out_tag_3; // @[STA_VDBB.scala 161:23:@12511.4 STA_VDBB.scala 181:29:@12674.4 STA_VDBB.scala 181:29:@12699.4 STA_VDBB.scala 181:29:@13466.4 STA_VDBB.scala 181:29:@13491.4 STA_VDBB.scala 181:29:@14258.4 STA_VDBB.scala 181:29:@14283.4 STA_VDBB.scala 181:29:@15050.4 STA_VDBB.scala 181:29:@15075.4 STA_VDBB.scala 181:29:@15842.4 STA_VDBB.scala 181:29:@15867.4 STA_VDBB.scala 181:29:@16634.4 STA_VDBB.scala 181:29:@16659.4 STA_VDBB.scala 181:29:@17426.4 STA_VDBB.scala 181:29:@17451.4 STA_VDBB.scala 181:29:@18218.4 STA_VDBB.scala 181:29:@18243.4 STA_VDBB.scala 293:23:@21343.4 STA_VDBB.scala 313:29:@21506.4 STA_VDBB.scala 313:29:@21531.4 STA_VDBB.scala 313:29:@22298.4 STA_VDBB.scala 313:29:@22323.4 STA_VDBB.scala 313:29:@23090.4 STA_VDBB.scala 313:29:@23115.4 STA_VDBB.scala 313:29:@23882.4 STA_VDBB.scala 313:29:@23907.4 STA_VDBB.scala 313:29:@24674.4 STA_VDBB.scala 313:29:@24699.4 STA_VDBB.scala 313:29:@25466.4 STA_VDBB.scala 313:29:@25491.4 STA_VDBB.scala 313:29:@26258.4 STA_VDBB.scala 313:29:@26283.4 STA_VDBB.scala 313:29:@27050.4 STA_VDBB.scala 313:29:@27075.4]
  assign ffb2_io_in_tag_1_4 = S8DP1_13_io_out_tag_4; // @[STA_VDBB.scala 161:23:@12512.4 STA_VDBB.scala 181:29:@12675.4 STA_VDBB.scala 181:29:@12700.4 STA_VDBB.scala 181:29:@13467.4 STA_VDBB.scala 181:29:@13492.4 STA_VDBB.scala 181:29:@14259.4 STA_VDBB.scala 181:29:@14284.4 STA_VDBB.scala 181:29:@15051.4 STA_VDBB.scala 181:29:@15076.4 STA_VDBB.scala 181:29:@15843.4 STA_VDBB.scala 181:29:@15868.4 STA_VDBB.scala 181:29:@16635.4 STA_VDBB.scala 181:29:@16660.4 STA_VDBB.scala 181:29:@17427.4 STA_VDBB.scala 181:29:@17452.4 STA_VDBB.scala 181:29:@18219.4 STA_VDBB.scala 181:29:@18244.4 STA_VDBB.scala 293:23:@21344.4 STA_VDBB.scala 313:29:@21507.4 STA_VDBB.scala 313:29:@21532.4 STA_VDBB.scala 313:29:@22299.4 STA_VDBB.scala 313:29:@22324.4 STA_VDBB.scala 313:29:@23091.4 STA_VDBB.scala 313:29:@23116.4 STA_VDBB.scala 313:29:@23883.4 STA_VDBB.scala 313:29:@23908.4 STA_VDBB.scala 313:29:@24675.4 STA_VDBB.scala 313:29:@24700.4 STA_VDBB.scala 313:29:@25467.4 STA_VDBB.scala 313:29:@25492.4 STA_VDBB.scala 313:29:@26259.4 STA_VDBB.scala 313:29:@26284.4 STA_VDBB.scala 313:29:@27051.4 STA_VDBB.scala 313:29:@27076.4]
  assign ffb2_io_in_tag_1_5 = S8DP1_13_io_out_tag_5; // @[STA_VDBB.scala 161:23:@12513.4 STA_VDBB.scala 181:29:@12676.4 STA_VDBB.scala 181:29:@12701.4 STA_VDBB.scala 181:29:@13468.4 STA_VDBB.scala 181:29:@13493.4 STA_VDBB.scala 181:29:@14260.4 STA_VDBB.scala 181:29:@14285.4 STA_VDBB.scala 181:29:@15052.4 STA_VDBB.scala 181:29:@15077.4 STA_VDBB.scala 181:29:@15844.4 STA_VDBB.scala 181:29:@15869.4 STA_VDBB.scala 181:29:@16636.4 STA_VDBB.scala 181:29:@16661.4 STA_VDBB.scala 181:29:@17428.4 STA_VDBB.scala 181:29:@17453.4 STA_VDBB.scala 181:29:@18220.4 STA_VDBB.scala 181:29:@18245.4 STA_VDBB.scala 293:23:@21345.4 STA_VDBB.scala 313:29:@21508.4 STA_VDBB.scala 313:29:@21533.4 STA_VDBB.scala 313:29:@22300.4 STA_VDBB.scala 313:29:@22325.4 STA_VDBB.scala 313:29:@23092.4 STA_VDBB.scala 313:29:@23117.4 STA_VDBB.scala 313:29:@23884.4 STA_VDBB.scala 313:29:@23909.4 STA_VDBB.scala 313:29:@24676.4 STA_VDBB.scala 313:29:@24701.4 STA_VDBB.scala 313:29:@25468.4 STA_VDBB.scala 313:29:@25493.4 STA_VDBB.scala 313:29:@26260.4 STA_VDBB.scala 313:29:@26285.4 STA_VDBB.scala 313:29:@27052.4 STA_VDBB.scala 313:29:@27077.4]
  assign ffb2_io_in_tag_1_6 = S8DP1_13_io_out_tag_6; // @[STA_VDBB.scala 161:23:@12514.4 STA_VDBB.scala 181:29:@12677.4 STA_VDBB.scala 181:29:@12702.4 STA_VDBB.scala 181:29:@13469.4 STA_VDBB.scala 181:29:@13494.4 STA_VDBB.scala 181:29:@14261.4 STA_VDBB.scala 181:29:@14286.4 STA_VDBB.scala 181:29:@15053.4 STA_VDBB.scala 181:29:@15078.4 STA_VDBB.scala 181:29:@15845.4 STA_VDBB.scala 181:29:@15870.4 STA_VDBB.scala 181:29:@16637.4 STA_VDBB.scala 181:29:@16662.4 STA_VDBB.scala 181:29:@17429.4 STA_VDBB.scala 181:29:@17454.4 STA_VDBB.scala 181:29:@18221.4 STA_VDBB.scala 181:29:@18246.4 STA_VDBB.scala 293:23:@21346.4 STA_VDBB.scala 313:29:@21509.4 STA_VDBB.scala 313:29:@21534.4 STA_VDBB.scala 313:29:@22301.4 STA_VDBB.scala 313:29:@22326.4 STA_VDBB.scala 313:29:@23093.4 STA_VDBB.scala 313:29:@23118.4 STA_VDBB.scala 313:29:@23885.4 STA_VDBB.scala 313:29:@23910.4 STA_VDBB.scala 313:29:@24677.4 STA_VDBB.scala 313:29:@24702.4 STA_VDBB.scala 313:29:@25469.4 STA_VDBB.scala 313:29:@25494.4 STA_VDBB.scala 313:29:@26261.4 STA_VDBB.scala 313:29:@26286.4 STA_VDBB.scala 313:29:@27053.4 STA_VDBB.scala 313:29:@27078.4]
  assign ffb2_io_in_tag_1_7 = S8DP1_13_io_out_tag_7; // @[STA_VDBB.scala 161:23:@12515.4 STA_VDBB.scala 181:29:@12678.4 STA_VDBB.scala 181:29:@12703.4 STA_VDBB.scala 181:29:@13470.4 STA_VDBB.scala 181:29:@13495.4 STA_VDBB.scala 181:29:@14262.4 STA_VDBB.scala 181:29:@14287.4 STA_VDBB.scala 181:29:@15054.4 STA_VDBB.scala 181:29:@15079.4 STA_VDBB.scala 181:29:@15846.4 STA_VDBB.scala 181:29:@15871.4 STA_VDBB.scala 181:29:@16638.4 STA_VDBB.scala 181:29:@16663.4 STA_VDBB.scala 181:29:@17430.4 STA_VDBB.scala 181:29:@17455.4 STA_VDBB.scala 181:29:@18222.4 STA_VDBB.scala 181:29:@18247.4 STA_VDBB.scala 293:23:@21347.4 STA_VDBB.scala 313:29:@21510.4 STA_VDBB.scala 313:29:@21535.4 STA_VDBB.scala 313:29:@22302.4 STA_VDBB.scala 313:29:@22327.4 STA_VDBB.scala 313:29:@23094.4 STA_VDBB.scala 313:29:@23119.4 STA_VDBB.scala 313:29:@23886.4 STA_VDBB.scala 313:29:@23911.4 STA_VDBB.scala 313:29:@24678.4 STA_VDBB.scala 313:29:@24703.4 STA_VDBB.scala 313:29:@25470.4 STA_VDBB.scala 313:29:@25495.4 STA_VDBB.scala 313:29:@26262.4 STA_VDBB.scala 313:29:@26287.4 STA_VDBB.scala 313:29:@27054.4 STA_VDBB.scala 313:29:@27079.4]
  assign ffb2_io_in_tag_2_0 = S8DP1_14_io_out_tag_0; // @[STA_VDBB.scala 161:23:@12532.4 STA_VDBB.scala 181:29:@12737.4 STA_VDBB.scala 181:29:@12762.4 STA_VDBB.scala 181:29:@13529.4 STA_VDBB.scala 181:29:@13554.4 STA_VDBB.scala 181:29:@14321.4 STA_VDBB.scala 181:29:@14346.4 STA_VDBB.scala 181:29:@15113.4 STA_VDBB.scala 181:29:@15138.4 STA_VDBB.scala 181:29:@15905.4 STA_VDBB.scala 181:29:@15930.4 STA_VDBB.scala 181:29:@16697.4 STA_VDBB.scala 181:29:@16722.4 STA_VDBB.scala 181:29:@17489.4 STA_VDBB.scala 181:29:@17514.4 STA_VDBB.scala 181:29:@18281.4 STA_VDBB.scala 181:29:@18306.4 STA_VDBB.scala 293:23:@21364.4 STA_VDBB.scala 313:29:@21569.4 STA_VDBB.scala 313:29:@21594.4 STA_VDBB.scala 313:29:@22361.4 STA_VDBB.scala 313:29:@22386.4 STA_VDBB.scala 313:29:@23153.4 STA_VDBB.scala 313:29:@23178.4 STA_VDBB.scala 313:29:@23945.4 STA_VDBB.scala 313:29:@23970.4 STA_VDBB.scala 313:29:@24737.4 STA_VDBB.scala 313:29:@24762.4 STA_VDBB.scala 313:29:@25529.4 STA_VDBB.scala 313:29:@25554.4 STA_VDBB.scala 313:29:@26321.4 STA_VDBB.scala 313:29:@26346.4 STA_VDBB.scala 313:29:@27113.4 STA_VDBB.scala 313:29:@27138.4]
  assign ffb2_io_in_tag_2_1 = S8DP1_14_io_out_tag_1; // @[STA_VDBB.scala 161:23:@12533.4 STA_VDBB.scala 181:29:@12738.4 STA_VDBB.scala 181:29:@12763.4 STA_VDBB.scala 181:29:@13530.4 STA_VDBB.scala 181:29:@13555.4 STA_VDBB.scala 181:29:@14322.4 STA_VDBB.scala 181:29:@14347.4 STA_VDBB.scala 181:29:@15114.4 STA_VDBB.scala 181:29:@15139.4 STA_VDBB.scala 181:29:@15906.4 STA_VDBB.scala 181:29:@15931.4 STA_VDBB.scala 181:29:@16698.4 STA_VDBB.scala 181:29:@16723.4 STA_VDBB.scala 181:29:@17490.4 STA_VDBB.scala 181:29:@17515.4 STA_VDBB.scala 181:29:@18282.4 STA_VDBB.scala 181:29:@18307.4 STA_VDBB.scala 293:23:@21365.4 STA_VDBB.scala 313:29:@21570.4 STA_VDBB.scala 313:29:@21595.4 STA_VDBB.scala 313:29:@22362.4 STA_VDBB.scala 313:29:@22387.4 STA_VDBB.scala 313:29:@23154.4 STA_VDBB.scala 313:29:@23179.4 STA_VDBB.scala 313:29:@23946.4 STA_VDBB.scala 313:29:@23971.4 STA_VDBB.scala 313:29:@24738.4 STA_VDBB.scala 313:29:@24763.4 STA_VDBB.scala 313:29:@25530.4 STA_VDBB.scala 313:29:@25555.4 STA_VDBB.scala 313:29:@26322.4 STA_VDBB.scala 313:29:@26347.4 STA_VDBB.scala 313:29:@27114.4 STA_VDBB.scala 313:29:@27139.4]
  assign ffb2_io_in_tag_2_2 = S8DP1_14_io_out_tag_2; // @[STA_VDBB.scala 161:23:@12534.4 STA_VDBB.scala 181:29:@12739.4 STA_VDBB.scala 181:29:@12764.4 STA_VDBB.scala 181:29:@13531.4 STA_VDBB.scala 181:29:@13556.4 STA_VDBB.scala 181:29:@14323.4 STA_VDBB.scala 181:29:@14348.4 STA_VDBB.scala 181:29:@15115.4 STA_VDBB.scala 181:29:@15140.4 STA_VDBB.scala 181:29:@15907.4 STA_VDBB.scala 181:29:@15932.4 STA_VDBB.scala 181:29:@16699.4 STA_VDBB.scala 181:29:@16724.4 STA_VDBB.scala 181:29:@17491.4 STA_VDBB.scala 181:29:@17516.4 STA_VDBB.scala 181:29:@18283.4 STA_VDBB.scala 181:29:@18308.4 STA_VDBB.scala 293:23:@21366.4 STA_VDBB.scala 313:29:@21571.4 STA_VDBB.scala 313:29:@21596.4 STA_VDBB.scala 313:29:@22363.4 STA_VDBB.scala 313:29:@22388.4 STA_VDBB.scala 313:29:@23155.4 STA_VDBB.scala 313:29:@23180.4 STA_VDBB.scala 313:29:@23947.4 STA_VDBB.scala 313:29:@23972.4 STA_VDBB.scala 313:29:@24739.4 STA_VDBB.scala 313:29:@24764.4 STA_VDBB.scala 313:29:@25531.4 STA_VDBB.scala 313:29:@25556.4 STA_VDBB.scala 313:29:@26323.4 STA_VDBB.scala 313:29:@26348.4 STA_VDBB.scala 313:29:@27115.4 STA_VDBB.scala 313:29:@27140.4]
  assign ffb2_io_in_tag_2_3 = S8DP1_14_io_out_tag_3; // @[STA_VDBB.scala 161:23:@12535.4 STA_VDBB.scala 181:29:@12740.4 STA_VDBB.scala 181:29:@12765.4 STA_VDBB.scala 181:29:@13532.4 STA_VDBB.scala 181:29:@13557.4 STA_VDBB.scala 181:29:@14324.4 STA_VDBB.scala 181:29:@14349.4 STA_VDBB.scala 181:29:@15116.4 STA_VDBB.scala 181:29:@15141.4 STA_VDBB.scala 181:29:@15908.4 STA_VDBB.scala 181:29:@15933.4 STA_VDBB.scala 181:29:@16700.4 STA_VDBB.scala 181:29:@16725.4 STA_VDBB.scala 181:29:@17492.4 STA_VDBB.scala 181:29:@17517.4 STA_VDBB.scala 181:29:@18284.4 STA_VDBB.scala 181:29:@18309.4 STA_VDBB.scala 293:23:@21367.4 STA_VDBB.scala 313:29:@21572.4 STA_VDBB.scala 313:29:@21597.4 STA_VDBB.scala 313:29:@22364.4 STA_VDBB.scala 313:29:@22389.4 STA_VDBB.scala 313:29:@23156.4 STA_VDBB.scala 313:29:@23181.4 STA_VDBB.scala 313:29:@23948.4 STA_VDBB.scala 313:29:@23973.4 STA_VDBB.scala 313:29:@24740.4 STA_VDBB.scala 313:29:@24765.4 STA_VDBB.scala 313:29:@25532.4 STA_VDBB.scala 313:29:@25557.4 STA_VDBB.scala 313:29:@26324.4 STA_VDBB.scala 313:29:@26349.4 STA_VDBB.scala 313:29:@27116.4 STA_VDBB.scala 313:29:@27141.4]
  assign ffb2_io_in_tag_2_4 = S8DP1_14_io_out_tag_4; // @[STA_VDBB.scala 161:23:@12536.4 STA_VDBB.scala 181:29:@12741.4 STA_VDBB.scala 181:29:@12766.4 STA_VDBB.scala 181:29:@13533.4 STA_VDBB.scala 181:29:@13558.4 STA_VDBB.scala 181:29:@14325.4 STA_VDBB.scala 181:29:@14350.4 STA_VDBB.scala 181:29:@15117.4 STA_VDBB.scala 181:29:@15142.4 STA_VDBB.scala 181:29:@15909.4 STA_VDBB.scala 181:29:@15934.4 STA_VDBB.scala 181:29:@16701.4 STA_VDBB.scala 181:29:@16726.4 STA_VDBB.scala 181:29:@17493.4 STA_VDBB.scala 181:29:@17518.4 STA_VDBB.scala 181:29:@18285.4 STA_VDBB.scala 181:29:@18310.4 STA_VDBB.scala 293:23:@21368.4 STA_VDBB.scala 313:29:@21573.4 STA_VDBB.scala 313:29:@21598.4 STA_VDBB.scala 313:29:@22365.4 STA_VDBB.scala 313:29:@22390.4 STA_VDBB.scala 313:29:@23157.4 STA_VDBB.scala 313:29:@23182.4 STA_VDBB.scala 313:29:@23949.4 STA_VDBB.scala 313:29:@23974.4 STA_VDBB.scala 313:29:@24741.4 STA_VDBB.scala 313:29:@24766.4 STA_VDBB.scala 313:29:@25533.4 STA_VDBB.scala 313:29:@25558.4 STA_VDBB.scala 313:29:@26325.4 STA_VDBB.scala 313:29:@26350.4 STA_VDBB.scala 313:29:@27117.4 STA_VDBB.scala 313:29:@27142.4]
  assign ffb2_io_in_tag_2_5 = S8DP1_14_io_out_tag_5; // @[STA_VDBB.scala 161:23:@12537.4 STA_VDBB.scala 181:29:@12742.4 STA_VDBB.scala 181:29:@12767.4 STA_VDBB.scala 181:29:@13534.4 STA_VDBB.scala 181:29:@13559.4 STA_VDBB.scala 181:29:@14326.4 STA_VDBB.scala 181:29:@14351.4 STA_VDBB.scala 181:29:@15118.4 STA_VDBB.scala 181:29:@15143.4 STA_VDBB.scala 181:29:@15910.4 STA_VDBB.scala 181:29:@15935.4 STA_VDBB.scala 181:29:@16702.4 STA_VDBB.scala 181:29:@16727.4 STA_VDBB.scala 181:29:@17494.4 STA_VDBB.scala 181:29:@17519.4 STA_VDBB.scala 181:29:@18286.4 STA_VDBB.scala 181:29:@18311.4 STA_VDBB.scala 293:23:@21369.4 STA_VDBB.scala 313:29:@21574.4 STA_VDBB.scala 313:29:@21599.4 STA_VDBB.scala 313:29:@22366.4 STA_VDBB.scala 313:29:@22391.4 STA_VDBB.scala 313:29:@23158.4 STA_VDBB.scala 313:29:@23183.4 STA_VDBB.scala 313:29:@23950.4 STA_VDBB.scala 313:29:@23975.4 STA_VDBB.scala 313:29:@24742.4 STA_VDBB.scala 313:29:@24767.4 STA_VDBB.scala 313:29:@25534.4 STA_VDBB.scala 313:29:@25559.4 STA_VDBB.scala 313:29:@26326.4 STA_VDBB.scala 313:29:@26351.4 STA_VDBB.scala 313:29:@27118.4 STA_VDBB.scala 313:29:@27143.4]
  assign ffb2_io_in_tag_2_6 = S8DP1_14_io_out_tag_6; // @[STA_VDBB.scala 161:23:@12538.4 STA_VDBB.scala 181:29:@12743.4 STA_VDBB.scala 181:29:@12768.4 STA_VDBB.scala 181:29:@13535.4 STA_VDBB.scala 181:29:@13560.4 STA_VDBB.scala 181:29:@14327.4 STA_VDBB.scala 181:29:@14352.4 STA_VDBB.scala 181:29:@15119.4 STA_VDBB.scala 181:29:@15144.4 STA_VDBB.scala 181:29:@15911.4 STA_VDBB.scala 181:29:@15936.4 STA_VDBB.scala 181:29:@16703.4 STA_VDBB.scala 181:29:@16728.4 STA_VDBB.scala 181:29:@17495.4 STA_VDBB.scala 181:29:@17520.4 STA_VDBB.scala 181:29:@18287.4 STA_VDBB.scala 181:29:@18312.4 STA_VDBB.scala 293:23:@21370.4 STA_VDBB.scala 313:29:@21575.4 STA_VDBB.scala 313:29:@21600.4 STA_VDBB.scala 313:29:@22367.4 STA_VDBB.scala 313:29:@22392.4 STA_VDBB.scala 313:29:@23159.4 STA_VDBB.scala 313:29:@23184.4 STA_VDBB.scala 313:29:@23951.4 STA_VDBB.scala 313:29:@23976.4 STA_VDBB.scala 313:29:@24743.4 STA_VDBB.scala 313:29:@24768.4 STA_VDBB.scala 313:29:@25535.4 STA_VDBB.scala 313:29:@25560.4 STA_VDBB.scala 313:29:@26327.4 STA_VDBB.scala 313:29:@26352.4 STA_VDBB.scala 313:29:@27119.4 STA_VDBB.scala 313:29:@27144.4]
  assign ffb2_io_in_tag_2_7 = S8DP1_14_io_out_tag_7; // @[STA_VDBB.scala 161:23:@12539.4 STA_VDBB.scala 181:29:@12744.4 STA_VDBB.scala 181:29:@12769.4 STA_VDBB.scala 181:29:@13536.4 STA_VDBB.scala 181:29:@13561.4 STA_VDBB.scala 181:29:@14328.4 STA_VDBB.scala 181:29:@14353.4 STA_VDBB.scala 181:29:@15120.4 STA_VDBB.scala 181:29:@15145.4 STA_VDBB.scala 181:29:@15912.4 STA_VDBB.scala 181:29:@15937.4 STA_VDBB.scala 181:29:@16704.4 STA_VDBB.scala 181:29:@16729.4 STA_VDBB.scala 181:29:@17496.4 STA_VDBB.scala 181:29:@17521.4 STA_VDBB.scala 181:29:@18288.4 STA_VDBB.scala 181:29:@18313.4 STA_VDBB.scala 293:23:@21371.4 STA_VDBB.scala 313:29:@21576.4 STA_VDBB.scala 313:29:@21601.4 STA_VDBB.scala 313:29:@22368.4 STA_VDBB.scala 313:29:@22393.4 STA_VDBB.scala 313:29:@23160.4 STA_VDBB.scala 313:29:@23185.4 STA_VDBB.scala 313:29:@23952.4 STA_VDBB.scala 313:29:@23977.4 STA_VDBB.scala 313:29:@24744.4 STA_VDBB.scala 313:29:@24769.4 STA_VDBB.scala 313:29:@25536.4 STA_VDBB.scala 313:29:@25561.4 STA_VDBB.scala 313:29:@26328.4 STA_VDBB.scala 313:29:@26353.4 STA_VDBB.scala 313:29:@27120.4 STA_VDBB.scala 313:29:@27145.4]
  assign ffb2_io_in_tag_3_0 = S8DP1_15_io_out_tag_0; // @[STA_VDBB.scala 161:23:@12556.4 STA_VDBB.scala 181:29:@12803.4 STA_VDBB.scala 181:29:@12828.4 STA_VDBB.scala 181:29:@13595.4 STA_VDBB.scala 181:29:@13620.4 STA_VDBB.scala 181:29:@14387.4 STA_VDBB.scala 181:29:@14412.4 STA_VDBB.scala 181:29:@15179.4 STA_VDBB.scala 181:29:@15204.4 STA_VDBB.scala 181:29:@15971.4 STA_VDBB.scala 181:29:@15996.4 STA_VDBB.scala 181:29:@16763.4 STA_VDBB.scala 181:29:@16788.4 STA_VDBB.scala 181:29:@17555.4 STA_VDBB.scala 181:29:@17580.4 STA_VDBB.scala 181:29:@18347.4 STA_VDBB.scala 181:29:@18372.4 STA_VDBB.scala 293:23:@21388.4 STA_VDBB.scala 313:29:@21635.4 STA_VDBB.scala 313:29:@21660.4 STA_VDBB.scala 313:29:@22427.4 STA_VDBB.scala 313:29:@22452.4 STA_VDBB.scala 313:29:@23219.4 STA_VDBB.scala 313:29:@23244.4 STA_VDBB.scala 313:29:@24011.4 STA_VDBB.scala 313:29:@24036.4 STA_VDBB.scala 313:29:@24803.4 STA_VDBB.scala 313:29:@24828.4 STA_VDBB.scala 313:29:@25595.4 STA_VDBB.scala 313:29:@25620.4 STA_VDBB.scala 313:29:@26387.4 STA_VDBB.scala 313:29:@26412.4 STA_VDBB.scala 313:29:@27179.4 STA_VDBB.scala 313:29:@27204.4]
  assign ffb2_io_in_tag_3_1 = S8DP1_15_io_out_tag_1; // @[STA_VDBB.scala 161:23:@12557.4 STA_VDBB.scala 181:29:@12804.4 STA_VDBB.scala 181:29:@12829.4 STA_VDBB.scala 181:29:@13596.4 STA_VDBB.scala 181:29:@13621.4 STA_VDBB.scala 181:29:@14388.4 STA_VDBB.scala 181:29:@14413.4 STA_VDBB.scala 181:29:@15180.4 STA_VDBB.scala 181:29:@15205.4 STA_VDBB.scala 181:29:@15972.4 STA_VDBB.scala 181:29:@15997.4 STA_VDBB.scala 181:29:@16764.4 STA_VDBB.scala 181:29:@16789.4 STA_VDBB.scala 181:29:@17556.4 STA_VDBB.scala 181:29:@17581.4 STA_VDBB.scala 181:29:@18348.4 STA_VDBB.scala 181:29:@18373.4 STA_VDBB.scala 293:23:@21389.4 STA_VDBB.scala 313:29:@21636.4 STA_VDBB.scala 313:29:@21661.4 STA_VDBB.scala 313:29:@22428.4 STA_VDBB.scala 313:29:@22453.4 STA_VDBB.scala 313:29:@23220.4 STA_VDBB.scala 313:29:@23245.4 STA_VDBB.scala 313:29:@24012.4 STA_VDBB.scala 313:29:@24037.4 STA_VDBB.scala 313:29:@24804.4 STA_VDBB.scala 313:29:@24829.4 STA_VDBB.scala 313:29:@25596.4 STA_VDBB.scala 313:29:@25621.4 STA_VDBB.scala 313:29:@26388.4 STA_VDBB.scala 313:29:@26413.4 STA_VDBB.scala 313:29:@27180.4 STA_VDBB.scala 313:29:@27205.4]
  assign ffb2_io_in_tag_3_2 = S8DP1_15_io_out_tag_2; // @[STA_VDBB.scala 161:23:@12558.4 STA_VDBB.scala 181:29:@12805.4 STA_VDBB.scala 181:29:@12830.4 STA_VDBB.scala 181:29:@13597.4 STA_VDBB.scala 181:29:@13622.4 STA_VDBB.scala 181:29:@14389.4 STA_VDBB.scala 181:29:@14414.4 STA_VDBB.scala 181:29:@15181.4 STA_VDBB.scala 181:29:@15206.4 STA_VDBB.scala 181:29:@15973.4 STA_VDBB.scala 181:29:@15998.4 STA_VDBB.scala 181:29:@16765.4 STA_VDBB.scala 181:29:@16790.4 STA_VDBB.scala 181:29:@17557.4 STA_VDBB.scala 181:29:@17582.4 STA_VDBB.scala 181:29:@18349.4 STA_VDBB.scala 181:29:@18374.4 STA_VDBB.scala 293:23:@21390.4 STA_VDBB.scala 313:29:@21637.4 STA_VDBB.scala 313:29:@21662.4 STA_VDBB.scala 313:29:@22429.4 STA_VDBB.scala 313:29:@22454.4 STA_VDBB.scala 313:29:@23221.4 STA_VDBB.scala 313:29:@23246.4 STA_VDBB.scala 313:29:@24013.4 STA_VDBB.scala 313:29:@24038.4 STA_VDBB.scala 313:29:@24805.4 STA_VDBB.scala 313:29:@24830.4 STA_VDBB.scala 313:29:@25597.4 STA_VDBB.scala 313:29:@25622.4 STA_VDBB.scala 313:29:@26389.4 STA_VDBB.scala 313:29:@26414.4 STA_VDBB.scala 313:29:@27181.4 STA_VDBB.scala 313:29:@27206.4]
  assign ffb2_io_in_tag_3_3 = S8DP1_15_io_out_tag_3; // @[STA_VDBB.scala 161:23:@12559.4 STA_VDBB.scala 181:29:@12806.4 STA_VDBB.scala 181:29:@12831.4 STA_VDBB.scala 181:29:@13598.4 STA_VDBB.scala 181:29:@13623.4 STA_VDBB.scala 181:29:@14390.4 STA_VDBB.scala 181:29:@14415.4 STA_VDBB.scala 181:29:@15182.4 STA_VDBB.scala 181:29:@15207.4 STA_VDBB.scala 181:29:@15974.4 STA_VDBB.scala 181:29:@15999.4 STA_VDBB.scala 181:29:@16766.4 STA_VDBB.scala 181:29:@16791.4 STA_VDBB.scala 181:29:@17558.4 STA_VDBB.scala 181:29:@17583.4 STA_VDBB.scala 181:29:@18350.4 STA_VDBB.scala 181:29:@18375.4 STA_VDBB.scala 293:23:@21391.4 STA_VDBB.scala 313:29:@21638.4 STA_VDBB.scala 313:29:@21663.4 STA_VDBB.scala 313:29:@22430.4 STA_VDBB.scala 313:29:@22455.4 STA_VDBB.scala 313:29:@23222.4 STA_VDBB.scala 313:29:@23247.4 STA_VDBB.scala 313:29:@24014.4 STA_VDBB.scala 313:29:@24039.4 STA_VDBB.scala 313:29:@24806.4 STA_VDBB.scala 313:29:@24831.4 STA_VDBB.scala 313:29:@25598.4 STA_VDBB.scala 313:29:@25623.4 STA_VDBB.scala 313:29:@26390.4 STA_VDBB.scala 313:29:@26415.4 STA_VDBB.scala 313:29:@27182.4 STA_VDBB.scala 313:29:@27207.4]
  assign ffb2_io_in_tag_3_4 = S8DP1_15_io_out_tag_4; // @[STA_VDBB.scala 161:23:@12560.4 STA_VDBB.scala 181:29:@12807.4 STA_VDBB.scala 181:29:@12832.4 STA_VDBB.scala 181:29:@13599.4 STA_VDBB.scala 181:29:@13624.4 STA_VDBB.scala 181:29:@14391.4 STA_VDBB.scala 181:29:@14416.4 STA_VDBB.scala 181:29:@15183.4 STA_VDBB.scala 181:29:@15208.4 STA_VDBB.scala 181:29:@15975.4 STA_VDBB.scala 181:29:@16000.4 STA_VDBB.scala 181:29:@16767.4 STA_VDBB.scala 181:29:@16792.4 STA_VDBB.scala 181:29:@17559.4 STA_VDBB.scala 181:29:@17584.4 STA_VDBB.scala 181:29:@18351.4 STA_VDBB.scala 181:29:@18376.4 STA_VDBB.scala 293:23:@21392.4 STA_VDBB.scala 313:29:@21639.4 STA_VDBB.scala 313:29:@21664.4 STA_VDBB.scala 313:29:@22431.4 STA_VDBB.scala 313:29:@22456.4 STA_VDBB.scala 313:29:@23223.4 STA_VDBB.scala 313:29:@23248.4 STA_VDBB.scala 313:29:@24015.4 STA_VDBB.scala 313:29:@24040.4 STA_VDBB.scala 313:29:@24807.4 STA_VDBB.scala 313:29:@24832.4 STA_VDBB.scala 313:29:@25599.4 STA_VDBB.scala 313:29:@25624.4 STA_VDBB.scala 313:29:@26391.4 STA_VDBB.scala 313:29:@26416.4 STA_VDBB.scala 313:29:@27183.4 STA_VDBB.scala 313:29:@27208.4]
  assign ffb2_io_in_tag_3_5 = S8DP1_15_io_out_tag_5; // @[STA_VDBB.scala 161:23:@12561.4 STA_VDBB.scala 181:29:@12808.4 STA_VDBB.scala 181:29:@12833.4 STA_VDBB.scala 181:29:@13600.4 STA_VDBB.scala 181:29:@13625.4 STA_VDBB.scala 181:29:@14392.4 STA_VDBB.scala 181:29:@14417.4 STA_VDBB.scala 181:29:@15184.4 STA_VDBB.scala 181:29:@15209.4 STA_VDBB.scala 181:29:@15976.4 STA_VDBB.scala 181:29:@16001.4 STA_VDBB.scala 181:29:@16768.4 STA_VDBB.scala 181:29:@16793.4 STA_VDBB.scala 181:29:@17560.4 STA_VDBB.scala 181:29:@17585.4 STA_VDBB.scala 181:29:@18352.4 STA_VDBB.scala 181:29:@18377.4 STA_VDBB.scala 293:23:@21393.4 STA_VDBB.scala 313:29:@21640.4 STA_VDBB.scala 313:29:@21665.4 STA_VDBB.scala 313:29:@22432.4 STA_VDBB.scala 313:29:@22457.4 STA_VDBB.scala 313:29:@23224.4 STA_VDBB.scala 313:29:@23249.4 STA_VDBB.scala 313:29:@24016.4 STA_VDBB.scala 313:29:@24041.4 STA_VDBB.scala 313:29:@24808.4 STA_VDBB.scala 313:29:@24833.4 STA_VDBB.scala 313:29:@25600.4 STA_VDBB.scala 313:29:@25625.4 STA_VDBB.scala 313:29:@26392.4 STA_VDBB.scala 313:29:@26417.4 STA_VDBB.scala 313:29:@27184.4 STA_VDBB.scala 313:29:@27209.4]
  assign ffb2_io_in_tag_3_6 = S8DP1_15_io_out_tag_6; // @[STA_VDBB.scala 161:23:@12562.4 STA_VDBB.scala 181:29:@12809.4 STA_VDBB.scala 181:29:@12834.4 STA_VDBB.scala 181:29:@13601.4 STA_VDBB.scala 181:29:@13626.4 STA_VDBB.scala 181:29:@14393.4 STA_VDBB.scala 181:29:@14418.4 STA_VDBB.scala 181:29:@15185.4 STA_VDBB.scala 181:29:@15210.4 STA_VDBB.scala 181:29:@15977.4 STA_VDBB.scala 181:29:@16002.4 STA_VDBB.scala 181:29:@16769.4 STA_VDBB.scala 181:29:@16794.4 STA_VDBB.scala 181:29:@17561.4 STA_VDBB.scala 181:29:@17586.4 STA_VDBB.scala 181:29:@18353.4 STA_VDBB.scala 181:29:@18378.4 STA_VDBB.scala 293:23:@21394.4 STA_VDBB.scala 313:29:@21641.4 STA_VDBB.scala 313:29:@21666.4 STA_VDBB.scala 313:29:@22433.4 STA_VDBB.scala 313:29:@22458.4 STA_VDBB.scala 313:29:@23225.4 STA_VDBB.scala 313:29:@23250.4 STA_VDBB.scala 313:29:@24017.4 STA_VDBB.scala 313:29:@24042.4 STA_VDBB.scala 313:29:@24809.4 STA_VDBB.scala 313:29:@24834.4 STA_VDBB.scala 313:29:@25601.4 STA_VDBB.scala 313:29:@25626.4 STA_VDBB.scala 313:29:@26393.4 STA_VDBB.scala 313:29:@26418.4 STA_VDBB.scala 313:29:@27185.4 STA_VDBB.scala 313:29:@27210.4]
  assign ffb2_io_in_tag_3_7 = S8DP1_15_io_out_tag_7; // @[STA_VDBB.scala 161:23:@12563.4 STA_VDBB.scala 181:29:@12810.4 STA_VDBB.scala 181:29:@12835.4 STA_VDBB.scala 181:29:@13602.4 STA_VDBB.scala 181:29:@13627.4 STA_VDBB.scala 181:29:@14394.4 STA_VDBB.scala 181:29:@14419.4 STA_VDBB.scala 181:29:@15186.4 STA_VDBB.scala 181:29:@15211.4 STA_VDBB.scala 181:29:@15978.4 STA_VDBB.scala 181:29:@16003.4 STA_VDBB.scala 181:29:@16770.4 STA_VDBB.scala 181:29:@16795.4 STA_VDBB.scala 181:29:@17562.4 STA_VDBB.scala 181:29:@17587.4 STA_VDBB.scala 181:29:@18354.4 STA_VDBB.scala 181:29:@18379.4 STA_VDBB.scala 293:23:@21395.4 STA_VDBB.scala 313:29:@21642.4 STA_VDBB.scala 313:29:@21667.4 STA_VDBB.scala 313:29:@22434.4 STA_VDBB.scala 313:29:@22459.4 STA_VDBB.scala 313:29:@23226.4 STA_VDBB.scala 313:29:@23251.4 STA_VDBB.scala 313:29:@24018.4 STA_VDBB.scala 313:29:@24043.4 STA_VDBB.scala 313:29:@24810.4 STA_VDBB.scala 313:29:@24835.4 STA_VDBB.scala 313:29:@25602.4 STA_VDBB.scala 313:29:@25627.4 STA_VDBB.scala 313:29:@26394.4 STA_VDBB.scala 313:29:@26419.4 STA_VDBB.scala 313:29:@27186.4 STA_VDBB.scala 313:29:@27211.4]
  assign ffa1_clock = clock; // @[:@9793.4]
  assign ffa1_reset = reset; // @[:@9794.4]
  assign ffa1_io_in_data_0_0 = io_in_A_0_8; // @[STA_VDBB.scala 92:29:@10076.4 STA_VDBB.scala 223:29:@18908.4]
  assign ffa1_io_in_data_0_1 = io_in_A_0_9; // @[STA_VDBB.scala 92:29:@10088.4 STA_VDBB.scala 223:29:@18920.4]
  assign ffa1_io_in_data_0_2 = io_in_A_0_10; // @[STA_VDBB.scala 92:29:@10100.4 STA_VDBB.scala 223:29:@18932.4]
  assign ffa1_io_in_data_0_3 = io_in_A_0_11; // @[STA_VDBB.scala 92:29:@10112.4 STA_VDBB.scala 223:29:@18944.4]
  assign ffa1_io_in_data_0_4 = io_in_A_0_12; // @[STA_VDBB.scala 92:29:@10124.4 STA_VDBB.scala 223:29:@18956.4]
  assign ffa1_io_in_data_0_5 = io_in_A_0_13; // @[STA_VDBB.scala 92:29:@10136.4 STA_VDBB.scala 223:29:@18968.4]
  assign ffa1_io_in_data_0_6 = io_in_A_0_14; // @[STA_VDBB.scala 92:29:@10148.4 STA_VDBB.scala 223:29:@18980.4]
  assign ffa1_io_in_data_0_7 = io_in_A_0_15; // @[STA_VDBB.scala 92:29:@10160.4 STA_VDBB.scala 223:29:@18992.4]
  assign ffa1_io_in_data_1_0 = io_in_A_1_8; // @[STA_VDBB.scala 92:29:@10078.4 STA_VDBB.scala 223:29:@18910.4]
  assign ffa1_io_in_data_1_1 = io_in_A_1_9; // @[STA_VDBB.scala 92:29:@10090.4 STA_VDBB.scala 223:29:@18922.4]
  assign ffa1_io_in_data_1_2 = io_in_A_1_10; // @[STA_VDBB.scala 92:29:@10102.4 STA_VDBB.scala 223:29:@18934.4]
  assign ffa1_io_in_data_1_3 = io_in_A_1_11; // @[STA_VDBB.scala 92:29:@10114.4 STA_VDBB.scala 223:29:@18946.4]
  assign ffa1_io_in_data_1_4 = io_in_A_1_12; // @[STA_VDBB.scala 92:29:@10126.4 STA_VDBB.scala 223:29:@18958.4]
  assign ffa1_io_in_data_1_5 = io_in_A_1_13; // @[STA_VDBB.scala 92:29:@10138.4 STA_VDBB.scala 223:29:@18970.4]
  assign ffa1_io_in_data_1_6 = io_in_A_1_14; // @[STA_VDBB.scala 92:29:@10150.4 STA_VDBB.scala 223:29:@18982.4]
  assign ffa1_io_in_data_1_7 = io_in_A_1_15; // @[STA_VDBB.scala 92:29:@10162.4 STA_VDBB.scala 223:29:@18994.4]
  assign ff00_clock = clock; // @[:@9796.4]
  assign ff00_reset = reset; // @[:@9797.4]
  assign ff00_io_in_data_0_0 = io_in_A_0_8; // @[STA_VDBB.scala 93:29:@10077.4 STA_VDBB.scala 224:29:@18909.4]
  assign ff00_io_in_data_0_1 = io_in_A_0_9; // @[STA_VDBB.scala 93:29:@10089.4 STA_VDBB.scala 224:29:@18921.4]
  assign ff00_io_in_data_0_2 = io_in_A_0_10; // @[STA_VDBB.scala 93:29:@10101.4 STA_VDBB.scala 224:29:@18933.4]
  assign ff00_io_in_data_0_3 = io_in_A_0_11; // @[STA_VDBB.scala 93:29:@10113.4 STA_VDBB.scala 224:29:@18945.4]
  assign ff00_io_in_data_0_4 = io_in_A_0_12; // @[STA_VDBB.scala 93:29:@10125.4 STA_VDBB.scala 224:29:@18957.4]
  assign ff00_io_in_data_0_5 = io_in_A_0_13; // @[STA_VDBB.scala 93:29:@10137.4 STA_VDBB.scala 224:29:@18969.4]
  assign ff00_io_in_data_0_6 = io_in_A_0_14; // @[STA_VDBB.scala 93:29:@10149.4 STA_VDBB.scala 224:29:@18981.4]
  assign ff00_io_in_data_0_7 = io_in_A_0_15; // @[STA_VDBB.scala 93:29:@10161.4 STA_VDBB.scala 224:29:@18993.4]
  assign ff00_io_in_data_1_0 = io_in_A_1_8; // @[STA_VDBB.scala 93:29:@10079.4 STA_VDBB.scala 224:29:@18911.4]
  assign ff00_io_in_data_1_1 = io_in_A_1_9; // @[STA_VDBB.scala 93:29:@10091.4 STA_VDBB.scala 224:29:@18923.4]
  assign ff00_io_in_data_1_2 = io_in_A_1_10; // @[STA_VDBB.scala 93:29:@10103.4 STA_VDBB.scala 224:29:@18935.4]
  assign ff00_io_in_data_1_3 = io_in_A_1_11; // @[STA_VDBB.scala 93:29:@10115.4 STA_VDBB.scala 224:29:@18947.4]
  assign ff00_io_in_data_1_4 = io_in_A_1_12; // @[STA_VDBB.scala 93:29:@10127.4 STA_VDBB.scala 224:29:@18959.4]
  assign ff00_io_in_data_1_5 = io_in_A_1_13; // @[STA_VDBB.scala 93:29:@10139.4 STA_VDBB.scala 224:29:@18971.4]
  assign ff00_io_in_data_1_6 = io_in_A_1_14; // @[STA_VDBB.scala 93:29:@10151.4 STA_VDBB.scala 224:29:@18983.4]
  assign ff00_io_in_data_1_7 = io_in_A_1_15; // @[STA_VDBB.scala 93:29:@10163.4 STA_VDBB.scala 224:29:@18995.4]
  assign ff01_clock = clock; // @[:@9799.4]
  assign ff01_reset = reset; // @[:@9800.4]
  assign ff01_io_in_data_0_0 = io_in_B_0_8; // @[STA_VDBB.scala 100:29:@10081.4 STA_VDBB.scala 234:29:@18913.4]
  assign ff01_io_in_data_0_1 = io_in_B_0_9; // @[STA_VDBB.scala 100:29:@10093.4 STA_VDBB.scala 234:29:@18925.4]
  assign ff01_io_in_data_0_2 = io_in_B_0_10; // @[STA_VDBB.scala 100:29:@10105.4 STA_VDBB.scala 234:29:@18937.4]
  assign ff01_io_in_data_0_3 = io_in_B_0_11; // @[STA_VDBB.scala 100:29:@10117.4 STA_VDBB.scala 234:29:@18949.4]
  assign ff01_io_in_data_0_4 = io_in_B_0_12; // @[STA_VDBB.scala 100:29:@10129.4 STA_VDBB.scala 234:29:@18961.4]
  assign ff01_io_in_data_0_5 = io_in_B_0_13; // @[STA_VDBB.scala 100:29:@10141.4 STA_VDBB.scala 234:29:@18973.4]
  assign ff01_io_in_data_0_6 = io_in_B_0_14; // @[STA_VDBB.scala 100:29:@10153.4 STA_VDBB.scala 234:29:@18985.4]
  assign ff01_io_in_data_0_7 = io_in_B_0_15; // @[STA_VDBB.scala 100:29:@10165.4 STA_VDBB.scala 234:29:@18997.4]
  assign ff01_io_in_data_1_0 = io_in_B_1_8; // @[STA_VDBB.scala 100:29:@10083.4 STA_VDBB.scala 234:29:@18915.4]
  assign ff01_io_in_data_1_1 = io_in_B_1_9; // @[STA_VDBB.scala 100:29:@10095.4 STA_VDBB.scala 234:29:@18927.4]
  assign ff01_io_in_data_1_2 = io_in_B_1_10; // @[STA_VDBB.scala 100:29:@10107.4 STA_VDBB.scala 234:29:@18939.4]
  assign ff01_io_in_data_1_3 = io_in_B_1_11; // @[STA_VDBB.scala 100:29:@10119.4 STA_VDBB.scala 234:29:@18951.4]
  assign ff01_io_in_data_1_4 = io_in_B_1_12; // @[STA_VDBB.scala 100:29:@10131.4 STA_VDBB.scala 234:29:@18963.4]
  assign ff01_io_in_data_1_5 = io_in_B_1_13; // @[STA_VDBB.scala 100:29:@10143.4 STA_VDBB.scala 234:29:@18975.4]
  assign ff01_io_in_data_1_6 = io_in_B_1_14; // @[STA_VDBB.scala 100:29:@10155.4 STA_VDBB.scala 234:29:@18987.4]
  assign ff01_io_in_data_1_7 = io_in_B_1_15; // @[STA_VDBB.scala 100:29:@10167.4 STA_VDBB.scala 234:29:@18999.4]
  assign ff01_io_in_data_2_0 = io_in_B_2_8; // @[STA_VDBB.scala 100:29:@10085.4 STA_VDBB.scala 234:29:@18917.4]
  assign ff01_io_in_data_2_1 = io_in_B_2_9; // @[STA_VDBB.scala 100:29:@10097.4 STA_VDBB.scala 234:29:@18929.4]
  assign ff01_io_in_data_2_2 = io_in_B_2_10; // @[STA_VDBB.scala 100:29:@10109.4 STA_VDBB.scala 234:29:@18941.4]
  assign ff01_io_in_data_2_3 = io_in_B_2_11; // @[STA_VDBB.scala 100:29:@10121.4 STA_VDBB.scala 234:29:@18953.4]
  assign ff01_io_in_data_2_4 = io_in_B_2_12; // @[STA_VDBB.scala 100:29:@10133.4 STA_VDBB.scala 234:29:@18965.4]
  assign ff01_io_in_data_2_5 = io_in_B_2_13; // @[STA_VDBB.scala 100:29:@10145.4 STA_VDBB.scala 234:29:@18977.4]
  assign ff01_io_in_data_2_6 = io_in_B_2_14; // @[STA_VDBB.scala 100:29:@10157.4 STA_VDBB.scala 234:29:@18989.4]
  assign ff01_io_in_data_2_7 = io_in_B_2_15; // @[STA_VDBB.scala 100:29:@10169.4 STA_VDBB.scala 234:29:@19001.4]
  assign ff01_io_in_data_3_0 = io_in_B_3_8; // @[STA_VDBB.scala 100:29:@10087.4 STA_VDBB.scala 234:29:@18919.4]
  assign ff01_io_in_data_3_1 = io_in_B_3_9; // @[STA_VDBB.scala 100:29:@10099.4 STA_VDBB.scala 234:29:@18931.4]
  assign ff01_io_in_data_3_2 = io_in_B_3_10; // @[STA_VDBB.scala 100:29:@10111.4 STA_VDBB.scala 234:29:@18943.4]
  assign ff01_io_in_data_3_3 = io_in_B_3_11; // @[STA_VDBB.scala 100:29:@10123.4 STA_VDBB.scala 234:29:@18955.4]
  assign ff01_io_in_data_3_4 = io_in_B_3_12; // @[STA_VDBB.scala 100:29:@10135.4 STA_VDBB.scala 234:29:@18967.4]
  assign ff01_io_in_data_3_5 = io_in_B_3_13; // @[STA_VDBB.scala 100:29:@10147.4 STA_VDBB.scala 234:29:@18979.4]
  assign ff01_io_in_data_3_6 = io_in_B_3_14; // @[STA_VDBB.scala 100:29:@10159.4 STA_VDBB.scala 234:29:@18991.4]
  assign ff01_io_in_data_3_7 = io_in_B_3_15; // @[STA_VDBB.scala 100:29:@10171.4 STA_VDBB.scala 234:29:@19003.4]
  assign ff01_io_in_tag_0_0 = S8DP1_24_io_out_tag_0; // @[STA_VDBB.scala 109:23:@10188.4 STA_VDBB.scala 194:29:@12869.4 STA_VDBB.scala 194:29:@12894.4 STA_VDBB.scala 194:29:@13661.4 STA_VDBB.scala 194:29:@13686.4 STA_VDBB.scala 194:29:@14453.4 STA_VDBB.scala 194:29:@14478.4 STA_VDBB.scala 194:29:@15245.4 STA_VDBB.scala 194:29:@15270.4 STA_VDBB.scala 194:29:@16037.4 STA_VDBB.scala 194:29:@16062.4 STA_VDBB.scala 194:29:@16829.4 STA_VDBB.scala 194:29:@16854.4 STA_VDBB.scala 194:29:@17621.4 STA_VDBB.scala 194:29:@17646.4 STA_VDBB.scala 194:29:@18413.4 STA_VDBB.scala 194:29:@18438.4 STA_VDBB.scala 242:23:@19020.4 STA_VDBB.scala 326:29:@21701.4 STA_VDBB.scala 326:29:@21726.4 STA_VDBB.scala 326:29:@22493.4 STA_VDBB.scala 326:29:@22518.4 STA_VDBB.scala 326:29:@23285.4 STA_VDBB.scala 326:29:@23310.4 STA_VDBB.scala 326:29:@24077.4 STA_VDBB.scala 326:29:@24102.4 STA_VDBB.scala 326:29:@24869.4 STA_VDBB.scala 326:29:@24894.4 STA_VDBB.scala 326:29:@25661.4 STA_VDBB.scala 326:29:@25686.4 STA_VDBB.scala 326:29:@26453.4 STA_VDBB.scala 326:29:@26478.4 STA_VDBB.scala 326:29:@27245.4 STA_VDBB.scala 326:29:@27270.4]
  assign ff01_io_in_tag_0_1 = S8DP1_24_io_out_tag_1; // @[STA_VDBB.scala 109:23:@10189.4 STA_VDBB.scala 194:29:@12870.4 STA_VDBB.scala 194:29:@12895.4 STA_VDBB.scala 194:29:@13662.4 STA_VDBB.scala 194:29:@13687.4 STA_VDBB.scala 194:29:@14454.4 STA_VDBB.scala 194:29:@14479.4 STA_VDBB.scala 194:29:@15246.4 STA_VDBB.scala 194:29:@15271.4 STA_VDBB.scala 194:29:@16038.4 STA_VDBB.scala 194:29:@16063.4 STA_VDBB.scala 194:29:@16830.4 STA_VDBB.scala 194:29:@16855.4 STA_VDBB.scala 194:29:@17622.4 STA_VDBB.scala 194:29:@17647.4 STA_VDBB.scala 194:29:@18414.4 STA_VDBB.scala 194:29:@18439.4 STA_VDBB.scala 242:23:@19021.4 STA_VDBB.scala 326:29:@21702.4 STA_VDBB.scala 326:29:@21727.4 STA_VDBB.scala 326:29:@22494.4 STA_VDBB.scala 326:29:@22519.4 STA_VDBB.scala 326:29:@23286.4 STA_VDBB.scala 326:29:@23311.4 STA_VDBB.scala 326:29:@24078.4 STA_VDBB.scala 326:29:@24103.4 STA_VDBB.scala 326:29:@24870.4 STA_VDBB.scala 326:29:@24895.4 STA_VDBB.scala 326:29:@25662.4 STA_VDBB.scala 326:29:@25687.4 STA_VDBB.scala 326:29:@26454.4 STA_VDBB.scala 326:29:@26479.4 STA_VDBB.scala 326:29:@27246.4 STA_VDBB.scala 326:29:@27271.4]
  assign ff01_io_in_tag_0_2 = S8DP1_24_io_out_tag_2; // @[STA_VDBB.scala 109:23:@10190.4 STA_VDBB.scala 194:29:@12871.4 STA_VDBB.scala 194:29:@12896.4 STA_VDBB.scala 194:29:@13663.4 STA_VDBB.scala 194:29:@13688.4 STA_VDBB.scala 194:29:@14455.4 STA_VDBB.scala 194:29:@14480.4 STA_VDBB.scala 194:29:@15247.4 STA_VDBB.scala 194:29:@15272.4 STA_VDBB.scala 194:29:@16039.4 STA_VDBB.scala 194:29:@16064.4 STA_VDBB.scala 194:29:@16831.4 STA_VDBB.scala 194:29:@16856.4 STA_VDBB.scala 194:29:@17623.4 STA_VDBB.scala 194:29:@17648.4 STA_VDBB.scala 194:29:@18415.4 STA_VDBB.scala 194:29:@18440.4 STA_VDBB.scala 242:23:@19022.4 STA_VDBB.scala 326:29:@21703.4 STA_VDBB.scala 326:29:@21728.4 STA_VDBB.scala 326:29:@22495.4 STA_VDBB.scala 326:29:@22520.4 STA_VDBB.scala 326:29:@23287.4 STA_VDBB.scala 326:29:@23312.4 STA_VDBB.scala 326:29:@24079.4 STA_VDBB.scala 326:29:@24104.4 STA_VDBB.scala 326:29:@24871.4 STA_VDBB.scala 326:29:@24896.4 STA_VDBB.scala 326:29:@25663.4 STA_VDBB.scala 326:29:@25688.4 STA_VDBB.scala 326:29:@26455.4 STA_VDBB.scala 326:29:@26480.4 STA_VDBB.scala 326:29:@27247.4 STA_VDBB.scala 326:29:@27272.4]
  assign ff01_io_in_tag_0_3 = S8DP1_24_io_out_tag_3; // @[STA_VDBB.scala 109:23:@10191.4 STA_VDBB.scala 194:29:@12872.4 STA_VDBB.scala 194:29:@12897.4 STA_VDBB.scala 194:29:@13664.4 STA_VDBB.scala 194:29:@13689.4 STA_VDBB.scala 194:29:@14456.4 STA_VDBB.scala 194:29:@14481.4 STA_VDBB.scala 194:29:@15248.4 STA_VDBB.scala 194:29:@15273.4 STA_VDBB.scala 194:29:@16040.4 STA_VDBB.scala 194:29:@16065.4 STA_VDBB.scala 194:29:@16832.4 STA_VDBB.scala 194:29:@16857.4 STA_VDBB.scala 194:29:@17624.4 STA_VDBB.scala 194:29:@17649.4 STA_VDBB.scala 194:29:@18416.4 STA_VDBB.scala 194:29:@18441.4 STA_VDBB.scala 242:23:@19023.4 STA_VDBB.scala 326:29:@21704.4 STA_VDBB.scala 326:29:@21729.4 STA_VDBB.scala 326:29:@22496.4 STA_VDBB.scala 326:29:@22521.4 STA_VDBB.scala 326:29:@23288.4 STA_VDBB.scala 326:29:@23313.4 STA_VDBB.scala 326:29:@24080.4 STA_VDBB.scala 326:29:@24105.4 STA_VDBB.scala 326:29:@24872.4 STA_VDBB.scala 326:29:@24897.4 STA_VDBB.scala 326:29:@25664.4 STA_VDBB.scala 326:29:@25689.4 STA_VDBB.scala 326:29:@26456.4 STA_VDBB.scala 326:29:@26481.4 STA_VDBB.scala 326:29:@27248.4 STA_VDBB.scala 326:29:@27273.4]
  assign ff01_io_in_tag_0_4 = S8DP1_24_io_out_tag_4; // @[STA_VDBB.scala 109:23:@10192.4 STA_VDBB.scala 194:29:@12873.4 STA_VDBB.scala 194:29:@12898.4 STA_VDBB.scala 194:29:@13665.4 STA_VDBB.scala 194:29:@13690.4 STA_VDBB.scala 194:29:@14457.4 STA_VDBB.scala 194:29:@14482.4 STA_VDBB.scala 194:29:@15249.4 STA_VDBB.scala 194:29:@15274.4 STA_VDBB.scala 194:29:@16041.4 STA_VDBB.scala 194:29:@16066.4 STA_VDBB.scala 194:29:@16833.4 STA_VDBB.scala 194:29:@16858.4 STA_VDBB.scala 194:29:@17625.4 STA_VDBB.scala 194:29:@17650.4 STA_VDBB.scala 194:29:@18417.4 STA_VDBB.scala 194:29:@18442.4 STA_VDBB.scala 242:23:@19024.4 STA_VDBB.scala 326:29:@21705.4 STA_VDBB.scala 326:29:@21730.4 STA_VDBB.scala 326:29:@22497.4 STA_VDBB.scala 326:29:@22522.4 STA_VDBB.scala 326:29:@23289.4 STA_VDBB.scala 326:29:@23314.4 STA_VDBB.scala 326:29:@24081.4 STA_VDBB.scala 326:29:@24106.4 STA_VDBB.scala 326:29:@24873.4 STA_VDBB.scala 326:29:@24898.4 STA_VDBB.scala 326:29:@25665.4 STA_VDBB.scala 326:29:@25690.4 STA_VDBB.scala 326:29:@26457.4 STA_VDBB.scala 326:29:@26482.4 STA_VDBB.scala 326:29:@27249.4 STA_VDBB.scala 326:29:@27274.4]
  assign ff01_io_in_tag_0_5 = S8DP1_24_io_out_tag_5; // @[STA_VDBB.scala 109:23:@10193.4 STA_VDBB.scala 194:29:@12874.4 STA_VDBB.scala 194:29:@12899.4 STA_VDBB.scala 194:29:@13666.4 STA_VDBB.scala 194:29:@13691.4 STA_VDBB.scala 194:29:@14458.4 STA_VDBB.scala 194:29:@14483.4 STA_VDBB.scala 194:29:@15250.4 STA_VDBB.scala 194:29:@15275.4 STA_VDBB.scala 194:29:@16042.4 STA_VDBB.scala 194:29:@16067.4 STA_VDBB.scala 194:29:@16834.4 STA_VDBB.scala 194:29:@16859.4 STA_VDBB.scala 194:29:@17626.4 STA_VDBB.scala 194:29:@17651.4 STA_VDBB.scala 194:29:@18418.4 STA_VDBB.scala 194:29:@18443.4 STA_VDBB.scala 242:23:@19025.4 STA_VDBB.scala 326:29:@21706.4 STA_VDBB.scala 326:29:@21731.4 STA_VDBB.scala 326:29:@22498.4 STA_VDBB.scala 326:29:@22523.4 STA_VDBB.scala 326:29:@23290.4 STA_VDBB.scala 326:29:@23315.4 STA_VDBB.scala 326:29:@24082.4 STA_VDBB.scala 326:29:@24107.4 STA_VDBB.scala 326:29:@24874.4 STA_VDBB.scala 326:29:@24899.4 STA_VDBB.scala 326:29:@25666.4 STA_VDBB.scala 326:29:@25691.4 STA_VDBB.scala 326:29:@26458.4 STA_VDBB.scala 326:29:@26483.4 STA_VDBB.scala 326:29:@27250.4 STA_VDBB.scala 326:29:@27275.4]
  assign ff01_io_in_tag_0_6 = S8DP1_24_io_out_tag_6; // @[STA_VDBB.scala 109:23:@10194.4 STA_VDBB.scala 194:29:@12875.4 STA_VDBB.scala 194:29:@12900.4 STA_VDBB.scala 194:29:@13667.4 STA_VDBB.scala 194:29:@13692.4 STA_VDBB.scala 194:29:@14459.4 STA_VDBB.scala 194:29:@14484.4 STA_VDBB.scala 194:29:@15251.4 STA_VDBB.scala 194:29:@15276.4 STA_VDBB.scala 194:29:@16043.4 STA_VDBB.scala 194:29:@16068.4 STA_VDBB.scala 194:29:@16835.4 STA_VDBB.scala 194:29:@16860.4 STA_VDBB.scala 194:29:@17627.4 STA_VDBB.scala 194:29:@17652.4 STA_VDBB.scala 194:29:@18419.4 STA_VDBB.scala 194:29:@18444.4 STA_VDBB.scala 242:23:@19026.4 STA_VDBB.scala 326:29:@21707.4 STA_VDBB.scala 326:29:@21732.4 STA_VDBB.scala 326:29:@22499.4 STA_VDBB.scala 326:29:@22524.4 STA_VDBB.scala 326:29:@23291.4 STA_VDBB.scala 326:29:@23316.4 STA_VDBB.scala 326:29:@24083.4 STA_VDBB.scala 326:29:@24108.4 STA_VDBB.scala 326:29:@24875.4 STA_VDBB.scala 326:29:@24900.4 STA_VDBB.scala 326:29:@25667.4 STA_VDBB.scala 326:29:@25692.4 STA_VDBB.scala 326:29:@26459.4 STA_VDBB.scala 326:29:@26484.4 STA_VDBB.scala 326:29:@27251.4 STA_VDBB.scala 326:29:@27276.4]
  assign ff01_io_in_tag_0_7 = S8DP1_24_io_out_tag_7; // @[STA_VDBB.scala 109:23:@10195.4 STA_VDBB.scala 194:29:@12876.4 STA_VDBB.scala 194:29:@12901.4 STA_VDBB.scala 194:29:@13668.4 STA_VDBB.scala 194:29:@13693.4 STA_VDBB.scala 194:29:@14460.4 STA_VDBB.scala 194:29:@14485.4 STA_VDBB.scala 194:29:@15252.4 STA_VDBB.scala 194:29:@15277.4 STA_VDBB.scala 194:29:@16044.4 STA_VDBB.scala 194:29:@16069.4 STA_VDBB.scala 194:29:@16836.4 STA_VDBB.scala 194:29:@16861.4 STA_VDBB.scala 194:29:@17628.4 STA_VDBB.scala 194:29:@17653.4 STA_VDBB.scala 194:29:@18420.4 STA_VDBB.scala 194:29:@18445.4 STA_VDBB.scala 242:23:@19027.4 STA_VDBB.scala 326:29:@21708.4 STA_VDBB.scala 326:29:@21733.4 STA_VDBB.scala 326:29:@22500.4 STA_VDBB.scala 326:29:@22525.4 STA_VDBB.scala 326:29:@23292.4 STA_VDBB.scala 326:29:@23317.4 STA_VDBB.scala 326:29:@24084.4 STA_VDBB.scala 326:29:@24109.4 STA_VDBB.scala 326:29:@24876.4 STA_VDBB.scala 326:29:@24901.4 STA_VDBB.scala 326:29:@25668.4 STA_VDBB.scala 326:29:@25693.4 STA_VDBB.scala 326:29:@26460.4 STA_VDBB.scala 326:29:@26485.4 STA_VDBB.scala 326:29:@27252.4 STA_VDBB.scala 326:29:@27277.4]
  assign ff01_io_in_tag_1_0 = S8DP1_25_io_out_tag_0; // @[STA_VDBB.scala 109:23:@10212.4 STA_VDBB.scala 194:29:@12935.4 STA_VDBB.scala 194:29:@12960.4 STA_VDBB.scala 194:29:@13727.4 STA_VDBB.scala 194:29:@13752.4 STA_VDBB.scala 194:29:@14519.4 STA_VDBB.scala 194:29:@14544.4 STA_VDBB.scala 194:29:@15311.4 STA_VDBB.scala 194:29:@15336.4 STA_VDBB.scala 194:29:@16103.4 STA_VDBB.scala 194:29:@16128.4 STA_VDBB.scala 194:29:@16895.4 STA_VDBB.scala 194:29:@16920.4 STA_VDBB.scala 194:29:@17687.4 STA_VDBB.scala 194:29:@17712.4 STA_VDBB.scala 194:29:@18479.4 STA_VDBB.scala 194:29:@18504.4 STA_VDBB.scala 242:23:@19044.4 STA_VDBB.scala 326:29:@21767.4 STA_VDBB.scala 326:29:@21792.4 STA_VDBB.scala 326:29:@22559.4 STA_VDBB.scala 326:29:@22584.4 STA_VDBB.scala 326:29:@23351.4 STA_VDBB.scala 326:29:@23376.4 STA_VDBB.scala 326:29:@24143.4 STA_VDBB.scala 326:29:@24168.4 STA_VDBB.scala 326:29:@24935.4 STA_VDBB.scala 326:29:@24960.4 STA_VDBB.scala 326:29:@25727.4 STA_VDBB.scala 326:29:@25752.4 STA_VDBB.scala 326:29:@26519.4 STA_VDBB.scala 326:29:@26544.4 STA_VDBB.scala 326:29:@27311.4 STA_VDBB.scala 326:29:@27336.4]
  assign ff01_io_in_tag_1_1 = S8DP1_25_io_out_tag_1; // @[STA_VDBB.scala 109:23:@10213.4 STA_VDBB.scala 194:29:@12936.4 STA_VDBB.scala 194:29:@12961.4 STA_VDBB.scala 194:29:@13728.4 STA_VDBB.scala 194:29:@13753.4 STA_VDBB.scala 194:29:@14520.4 STA_VDBB.scala 194:29:@14545.4 STA_VDBB.scala 194:29:@15312.4 STA_VDBB.scala 194:29:@15337.4 STA_VDBB.scala 194:29:@16104.4 STA_VDBB.scala 194:29:@16129.4 STA_VDBB.scala 194:29:@16896.4 STA_VDBB.scala 194:29:@16921.4 STA_VDBB.scala 194:29:@17688.4 STA_VDBB.scala 194:29:@17713.4 STA_VDBB.scala 194:29:@18480.4 STA_VDBB.scala 194:29:@18505.4 STA_VDBB.scala 242:23:@19045.4 STA_VDBB.scala 326:29:@21768.4 STA_VDBB.scala 326:29:@21793.4 STA_VDBB.scala 326:29:@22560.4 STA_VDBB.scala 326:29:@22585.4 STA_VDBB.scala 326:29:@23352.4 STA_VDBB.scala 326:29:@23377.4 STA_VDBB.scala 326:29:@24144.4 STA_VDBB.scala 326:29:@24169.4 STA_VDBB.scala 326:29:@24936.4 STA_VDBB.scala 326:29:@24961.4 STA_VDBB.scala 326:29:@25728.4 STA_VDBB.scala 326:29:@25753.4 STA_VDBB.scala 326:29:@26520.4 STA_VDBB.scala 326:29:@26545.4 STA_VDBB.scala 326:29:@27312.4 STA_VDBB.scala 326:29:@27337.4]
  assign ff01_io_in_tag_1_2 = S8DP1_25_io_out_tag_2; // @[STA_VDBB.scala 109:23:@10214.4 STA_VDBB.scala 194:29:@12937.4 STA_VDBB.scala 194:29:@12962.4 STA_VDBB.scala 194:29:@13729.4 STA_VDBB.scala 194:29:@13754.4 STA_VDBB.scala 194:29:@14521.4 STA_VDBB.scala 194:29:@14546.4 STA_VDBB.scala 194:29:@15313.4 STA_VDBB.scala 194:29:@15338.4 STA_VDBB.scala 194:29:@16105.4 STA_VDBB.scala 194:29:@16130.4 STA_VDBB.scala 194:29:@16897.4 STA_VDBB.scala 194:29:@16922.4 STA_VDBB.scala 194:29:@17689.4 STA_VDBB.scala 194:29:@17714.4 STA_VDBB.scala 194:29:@18481.4 STA_VDBB.scala 194:29:@18506.4 STA_VDBB.scala 242:23:@19046.4 STA_VDBB.scala 326:29:@21769.4 STA_VDBB.scala 326:29:@21794.4 STA_VDBB.scala 326:29:@22561.4 STA_VDBB.scala 326:29:@22586.4 STA_VDBB.scala 326:29:@23353.4 STA_VDBB.scala 326:29:@23378.4 STA_VDBB.scala 326:29:@24145.4 STA_VDBB.scala 326:29:@24170.4 STA_VDBB.scala 326:29:@24937.4 STA_VDBB.scala 326:29:@24962.4 STA_VDBB.scala 326:29:@25729.4 STA_VDBB.scala 326:29:@25754.4 STA_VDBB.scala 326:29:@26521.4 STA_VDBB.scala 326:29:@26546.4 STA_VDBB.scala 326:29:@27313.4 STA_VDBB.scala 326:29:@27338.4]
  assign ff01_io_in_tag_1_3 = S8DP1_25_io_out_tag_3; // @[STA_VDBB.scala 109:23:@10215.4 STA_VDBB.scala 194:29:@12938.4 STA_VDBB.scala 194:29:@12963.4 STA_VDBB.scala 194:29:@13730.4 STA_VDBB.scala 194:29:@13755.4 STA_VDBB.scala 194:29:@14522.4 STA_VDBB.scala 194:29:@14547.4 STA_VDBB.scala 194:29:@15314.4 STA_VDBB.scala 194:29:@15339.4 STA_VDBB.scala 194:29:@16106.4 STA_VDBB.scala 194:29:@16131.4 STA_VDBB.scala 194:29:@16898.4 STA_VDBB.scala 194:29:@16923.4 STA_VDBB.scala 194:29:@17690.4 STA_VDBB.scala 194:29:@17715.4 STA_VDBB.scala 194:29:@18482.4 STA_VDBB.scala 194:29:@18507.4 STA_VDBB.scala 242:23:@19047.4 STA_VDBB.scala 326:29:@21770.4 STA_VDBB.scala 326:29:@21795.4 STA_VDBB.scala 326:29:@22562.4 STA_VDBB.scala 326:29:@22587.4 STA_VDBB.scala 326:29:@23354.4 STA_VDBB.scala 326:29:@23379.4 STA_VDBB.scala 326:29:@24146.4 STA_VDBB.scala 326:29:@24171.4 STA_VDBB.scala 326:29:@24938.4 STA_VDBB.scala 326:29:@24963.4 STA_VDBB.scala 326:29:@25730.4 STA_VDBB.scala 326:29:@25755.4 STA_VDBB.scala 326:29:@26522.4 STA_VDBB.scala 326:29:@26547.4 STA_VDBB.scala 326:29:@27314.4 STA_VDBB.scala 326:29:@27339.4]
  assign ff01_io_in_tag_1_4 = S8DP1_25_io_out_tag_4; // @[STA_VDBB.scala 109:23:@10216.4 STA_VDBB.scala 194:29:@12939.4 STA_VDBB.scala 194:29:@12964.4 STA_VDBB.scala 194:29:@13731.4 STA_VDBB.scala 194:29:@13756.4 STA_VDBB.scala 194:29:@14523.4 STA_VDBB.scala 194:29:@14548.4 STA_VDBB.scala 194:29:@15315.4 STA_VDBB.scala 194:29:@15340.4 STA_VDBB.scala 194:29:@16107.4 STA_VDBB.scala 194:29:@16132.4 STA_VDBB.scala 194:29:@16899.4 STA_VDBB.scala 194:29:@16924.4 STA_VDBB.scala 194:29:@17691.4 STA_VDBB.scala 194:29:@17716.4 STA_VDBB.scala 194:29:@18483.4 STA_VDBB.scala 194:29:@18508.4 STA_VDBB.scala 242:23:@19048.4 STA_VDBB.scala 326:29:@21771.4 STA_VDBB.scala 326:29:@21796.4 STA_VDBB.scala 326:29:@22563.4 STA_VDBB.scala 326:29:@22588.4 STA_VDBB.scala 326:29:@23355.4 STA_VDBB.scala 326:29:@23380.4 STA_VDBB.scala 326:29:@24147.4 STA_VDBB.scala 326:29:@24172.4 STA_VDBB.scala 326:29:@24939.4 STA_VDBB.scala 326:29:@24964.4 STA_VDBB.scala 326:29:@25731.4 STA_VDBB.scala 326:29:@25756.4 STA_VDBB.scala 326:29:@26523.4 STA_VDBB.scala 326:29:@26548.4 STA_VDBB.scala 326:29:@27315.4 STA_VDBB.scala 326:29:@27340.4]
  assign ff01_io_in_tag_1_5 = S8DP1_25_io_out_tag_5; // @[STA_VDBB.scala 109:23:@10217.4 STA_VDBB.scala 194:29:@12940.4 STA_VDBB.scala 194:29:@12965.4 STA_VDBB.scala 194:29:@13732.4 STA_VDBB.scala 194:29:@13757.4 STA_VDBB.scala 194:29:@14524.4 STA_VDBB.scala 194:29:@14549.4 STA_VDBB.scala 194:29:@15316.4 STA_VDBB.scala 194:29:@15341.4 STA_VDBB.scala 194:29:@16108.4 STA_VDBB.scala 194:29:@16133.4 STA_VDBB.scala 194:29:@16900.4 STA_VDBB.scala 194:29:@16925.4 STA_VDBB.scala 194:29:@17692.4 STA_VDBB.scala 194:29:@17717.4 STA_VDBB.scala 194:29:@18484.4 STA_VDBB.scala 194:29:@18509.4 STA_VDBB.scala 242:23:@19049.4 STA_VDBB.scala 326:29:@21772.4 STA_VDBB.scala 326:29:@21797.4 STA_VDBB.scala 326:29:@22564.4 STA_VDBB.scala 326:29:@22589.4 STA_VDBB.scala 326:29:@23356.4 STA_VDBB.scala 326:29:@23381.4 STA_VDBB.scala 326:29:@24148.4 STA_VDBB.scala 326:29:@24173.4 STA_VDBB.scala 326:29:@24940.4 STA_VDBB.scala 326:29:@24965.4 STA_VDBB.scala 326:29:@25732.4 STA_VDBB.scala 326:29:@25757.4 STA_VDBB.scala 326:29:@26524.4 STA_VDBB.scala 326:29:@26549.4 STA_VDBB.scala 326:29:@27316.4 STA_VDBB.scala 326:29:@27341.4]
  assign ff01_io_in_tag_1_6 = S8DP1_25_io_out_tag_6; // @[STA_VDBB.scala 109:23:@10218.4 STA_VDBB.scala 194:29:@12941.4 STA_VDBB.scala 194:29:@12966.4 STA_VDBB.scala 194:29:@13733.4 STA_VDBB.scala 194:29:@13758.4 STA_VDBB.scala 194:29:@14525.4 STA_VDBB.scala 194:29:@14550.4 STA_VDBB.scala 194:29:@15317.4 STA_VDBB.scala 194:29:@15342.4 STA_VDBB.scala 194:29:@16109.4 STA_VDBB.scala 194:29:@16134.4 STA_VDBB.scala 194:29:@16901.4 STA_VDBB.scala 194:29:@16926.4 STA_VDBB.scala 194:29:@17693.4 STA_VDBB.scala 194:29:@17718.4 STA_VDBB.scala 194:29:@18485.4 STA_VDBB.scala 194:29:@18510.4 STA_VDBB.scala 242:23:@19050.4 STA_VDBB.scala 326:29:@21773.4 STA_VDBB.scala 326:29:@21798.4 STA_VDBB.scala 326:29:@22565.4 STA_VDBB.scala 326:29:@22590.4 STA_VDBB.scala 326:29:@23357.4 STA_VDBB.scala 326:29:@23382.4 STA_VDBB.scala 326:29:@24149.4 STA_VDBB.scala 326:29:@24174.4 STA_VDBB.scala 326:29:@24941.4 STA_VDBB.scala 326:29:@24966.4 STA_VDBB.scala 326:29:@25733.4 STA_VDBB.scala 326:29:@25758.4 STA_VDBB.scala 326:29:@26525.4 STA_VDBB.scala 326:29:@26550.4 STA_VDBB.scala 326:29:@27317.4 STA_VDBB.scala 326:29:@27342.4]
  assign ff01_io_in_tag_1_7 = S8DP1_25_io_out_tag_7; // @[STA_VDBB.scala 109:23:@10219.4 STA_VDBB.scala 194:29:@12942.4 STA_VDBB.scala 194:29:@12967.4 STA_VDBB.scala 194:29:@13734.4 STA_VDBB.scala 194:29:@13759.4 STA_VDBB.scala 194:29:@14526.4 STA_VDBB.scala 194:29:@14551.4 STA_VDBB.scala 194:29:@15318.4 STA_VDBB.scala 194:29:@15343.4 STA_VDBB.scala 194:29:@16110.4 STA_VDBB.scala 194:29:@16135.4 STA_VDBB.scala 194:29:@16902.4 STA_VDBB.scala 194:29:@16927.4 STA_VDBB.scala 194:29:@17694.4 STA_VDBB.scala 194:29:@17719.4 STA_VDBB.scala 194:29:@18486.4 STA_VDBB.scala 194:29:@18511.4 STA_VDBB.scala 242:23:@19051.4 STA_VDBB.scala 326:29:@21774.4 STA_VDBB.scala 326:29:@21799.4 STA_VDBB.scala 326:29:@22566.4 STA_VDBB.scala 326:29:@22591.4 STA_VDBB.scala 326:29:@23358.4 STA_VDBB.scala 326:29:@23383.4 STA_VDBB.scala 326:29:@24150.4 STA_VDBB.scala 326:29:@24175.4 STA_VDBB.scala 326:29:@24942.4 STA_VDBB.scala 326:29:@24967.4 STA_VDBB.scala 326:29:@25734.4 STA_VDBB.scala 326:29:@25759.4 STA_VDBB.scala 326:29:@26526.4 STA_VDBB.scala 326:29:@26551.4 STA_VDBB.scala 326:29:@27318.4 STA_VDBB.scala 326:29:@27343.4]
  assign ff01_io_in_tag_2_0 = S8DP1_26_io_out_tag_0; // @[STA_VDBB.scala 109:23:@10236.4 STA_VDBB.scala 194:29:@13001.4 STA_VDBB.scala 194:29:@13026.4 STA_VDBB.scala 194:29:@13793.4 STA_VDBB.scala 194:29:@13818.4 STA_VDBB.scala 194:29:@14585.4 STA_VDBB.scala 194:29:@14610.4 STA_VDBB.scala 194:29:@15377.4 STA_VDBB.scala 194:29:@15402.4 STA_VDBB.scala 194:29:@16169.4 STA_VDBB.scala 194:29:@16194.4 STA_VDBB.scala 194:29:@16961.4 STA_VDBB.scala 194:29:@16986.4 STA_VDBB.scala 194:29:@17753.4 STA_VDBB.scala 194:29:@17778.4 STA_VDBB.scala 194:29:@18545.4 STA_VDBB.scala 194:29:@18570.4 STA_VDBB.scala 242:23:@19068.4 STA_VDBB.scala 326:29:@21833.4 STA_VDBB.scala 326:29:@21858.4 STA_VDBB.scala 326:29:@22625.4 STA_VDBB.scala 326:29:@22650.4 STA_VDBB.scala 326:29:@23417.4 STA_VDBB.scala 326:29:@23442.4 STA_VDBB.scala 326:29:@24209.4 STA_VDBB.scala 326:29:@24234.4 STA_VDBB.scala 326:29:@25001.4 STA_VDBB.scala 326:29:@25026.4 STA_VDBB.scala 326:29:@25793.4 STA_VDBB.scala 326:29:@25818.4 STA_VDBB.scala 326:29:@26585.4 STA_VDBB.scala 326:29:@26610.4 STA_VDBB.scala 326:29:@27377.4 STA_VDBB.scala 326:29:@27402.4]
  assign ff01_io_in_tag_2_1 = S8DP1_26_io_out_tag_1; // @[STA_VDBB.scala 109:23:@10237.4 STA_VDBB.scala 194:29:@13002.4 STA_VDBB.scala 194:29:@13027.4 STA_VDBB.scala 194:29:@13794.4 STA_VDBB.scala 194:29:@13819.4 STA_VDBB.scala 194:29:@14586.4 STA_VDBB.scala 194:29:@14611.4 STA_VDBB.scala 194:29:@15378.4 STA_VDBB.scala 194:29:@15403.4 STA_VDBB.scala 194:29:@16170.4 STA_VDBB.scala 194:29:@16195.4 STA_VDBB.scala 194:29:@16962.4 STA_VDBB.scala 194:29:@16987.4 STA_VDBB.scala 194:29:@17754.4 STA_VDBB.scala 194:29:@17779.4 STA_VDBB.scala 194:29:@18546.4 STA_VDBB.scala 194:29:@18571.4 STA_VDBB.scala 242:23:@19069.4 STA_VDBB.scala 326:29:@21834.4 STA_VDBB.scala 326:29:@21859.4 STA_VDBB.scala 326:29:@22626.4 STA_VDBB.scala 326:29:@22651.4 STA_VDBB.scala 326:29:@23418.4 STA_VDBB.scala 326:29:@23443.4 STA_VDBB.scala 326:29:@24210.4 STA_VDBB.scala 326:29:@24235.4 STA_VDBB.scala 326:29:@25002.4 STA_VDBB.scala 326:29:@25027.4 STA_VDBB.scala 326:29:@25794.4 STA_VDBB.scala 326:29:@25819.4 STA_VDBB.scala 326:29:@26586.4 STA_VDBB.scala 326:29:@26611.4 STA_VDBB.scala 326:29:@27378.4 STA_VDBB.scala 326:29:@27403.4]
  assign ff01_io_in_tag_2_2 = S8DP1_26_io_out_tag_2; // @[STA_VDBB.scala 109:23:@10238.4 STA_VDBB.scala 194:29:@13003.4 STA_VDBB.scala 194:29:@13028.4 STA_VDBB.scala 194:29:@13795.4 STA_VDBB.scala 194:29:@13820.4 STA_VDBB.scala 194:29:@14587.4 STA_VDBB.scala 194:29:@14612.4 STA_VDBB.scala 194:29:@15379.4 STA_VDBB.scala 194:29:@15404.4 STA_VDBB.scala 194:29:@16171.4 STA_VDBB.scala 194:29:@16196.4 STA_VDBB.scala 194:29:@16963.4 STA_VDBB.scala 194:29:@16988.4 STA_VDBB.scala 194:29:@17755.4 STA_VDBB.scala 194:29:@17780.4 STA_VDBB.scala 194:29:@18547.4 STA_VDBB.scala 194:29:@18572.4 STA_VDBB.scala 242:23:@19070.4 STA_VDBB.scala 326:29:@21835.4 STA_VDBB.scala 326:29:@21860.4 STA_VDBB.scala 326:29:@22627.4 STA_VDBB.scala 326:29:@22652.4 STA_VDBB.scala 326:29:@23419.4 STA_VDBB.scala 326:29:@23444.4 STA_VDBB.scala 326:29:@24211.4 STA_VDBB.scala 326:29:@24236.4 STA_VDBB.scala 326:29:@25003.4 STA_VDBB.scala 326:29:@25028.4 STA_VDBB.scala 326:29:@25795.4 STA_VDBB.scala 326:29:@25820.4 STA_VDBB.scala 326:29:@26587.4 STA_VDBB.scala 326:29:@26612.4 STA_VDBB.scala 326:29:@27379.4 STA_VDBB.scala 326:29:@27404.4]
  assign ff01_io_in_tag_2_3 = S8DP1_26_io_out_tag_3; // @[STA_VDBB.scala 109:23:@10239.4 STA_VDBB.scala 194:29:@13004.4 STA_VDBB.scala 194:29:@13029.4 STA_VDBB.scala 194:29:@13796.4 STA_VDBB.scala 194:29:@13821.4 STA_VDBB.scala 194:29:@14588.4 STA_VDBB.scala 194:29:@14613.4 STA_VDBB.scala 194:29:@15380.4 STA_VDBB.scala 194:29:@15405.4 STA_VDBB.scala 194:29:@16172.4 STA_VDBB.scala 194:29:@16197.4 STA_VDBB.scala 194:29:@16964.4 STA_VDBB.scala 194:29:@16989.4 STA_VDBB.scala 194:29:@17756.4 STA_VDBB.scala 194:29:@17781.4 STA_VDBB.scala 194:29:@18548.4 STA_VDBB.scala 194:29:@18573.4 STA_VDBB.scala 242:23:@19071.4 STA_VDBB.scala 326:29:@21836.4 STA_VDBB.scala 326:29:@21861.4 STA_VDBB.scala 326:29:@22628.4 STA_VDBB.scala 326:29:@22653.4 STA_VDBB.scala 326:29:@23420.4 STA_VDBB.scala 326:29:@23445.4 STA_VDBB.scala 326:29:@24212.4 STA_VDBB.scala 326:29:@24237.4 STA_VDBB.scala 326:29:@25004.4 STA_VDBB.scala 326:29:@25029.4 STA_VDBB.scala 326:29:@25796.4 STA_VDBB.scala 326:29:@25821.4 STA_VDBB.scala 326:29:@26588.4 STA_VDBB.scala 326:29:@26613.4 STA_VDBB.scala 326:29:@27380.4 STA_VDBB.scala 326:29:@27405.4]
  assign ff01_io_in_tag_2_4 = S8DP1_26_io_out_tag_4; // @[STA_VDBB.scala 109:23:@10240.4 STA_VDBB.scala 194:29:@13005.4 STA_VDBB.scala 194:29:@13030.4 STA_VDBB.scala 194:29:@13797.4 STA_VDBB.scala 194:29:@13822.4 STA_VDBB.scala 194:29:@14589.4 STA_VDBB.scala 194:29:@14614.4 STA_VDBB.scala 194:29:@15381.4 STA_VDBB.scala 194:29:@15406.4 STA_VDBB.scala 194:29:@16173.4 STA_VDBB.scala 194:29:@16198.4 STA_VDBB.scala 194:29:@16965.4 STA_VDBB.scala 194:29:@16990.4 STA_VDBB.scala 194:29:@17757.4 STA_VDBB.scala 194:29:@17782.4 STA_VDBB.scala 194:29:@18549.4 STA_VDBB.scala 194:29:@18574.4 STA_VDBB.scala 242:23:@19072.4 STA_VDBB.scala 326:29:@21837.4 STA_VDBB.scala 326:29:@21862.4 STA_VDBB.scala 326:29:@22629.4 STA_VDBB.scala 326:29:@22654.4 STA_VDBB.scala 326:29:@23421.4 STA_VDBB.scala 326:29:@23446.4 STA_VDBB.scala 326:29:@24213.4 STA_VDBB.scala 326:29:@24238.4 STA_VDBB.scala 326:29:@25005.4 STA_VDBB.scala 326:29:@25030.4 STA_VDBB.scala 326:29:@25797.4 STA_VDBB.scala 326:29:@25822.4 STA_VDBB.scala 326:29:@26589.4 STA_VDBB.scala 326:29:@26614.4 STA_VDBB.scala 326:29:@27381.4 STA_VDBB.scala 326:29:@27406.4]
  assign ff01_io_in_tag_2_5 = S8DP1_26_io_out_tag_5; // @[STA_VDBB.scala 109:23:@10241.4 STA_VDBB.scala 194:29:@13006.4 STA_VDBB.scala 194:29:@13031.4 STA_VDBB.scala 194:29:@13798.4 STA_VDBB.scala 194:29:@13823.4 STA_VDBB.scala 194:29:@14590.4 STA_VDBB.scala 194:29:@14615.4 STA_VDBB.scala 194:29:@15382.4 STA_VDBB.scala 194:29:@15407.4 STA_VDBB.scala 194:29:@16174.4 STA_VDBB.scala 194:29:@16199.4 STA_VDBB.scala 194:29:@16966.4 STA_VDBB.scala 194:29:@16991.4 STA_VDBB.scala 194:29:@17758.4 STA_VDBB.scala 194:29:@17783.4 STA_VDBB.scala 194:29:@18550.4 STA_VDBB.scala 194:29:@18575.4 STA_VDBB.scala 242:23:@19073.4 STA_VDBB.scala 326:29:@21838.4 STA_VDBB.scala 326:29:@21863.4 STA_VDBB.scala 326:29:@22630.4 STA_VDBB.scala 326:29:@22655.4 STA_VDBB.scala 326:29:@23422.4 STA_VDBB.scala 326:29:@23447.4 STA_VDBB.scala 326:29:@24214.4 STA_VDBB.scala 326:29:@24239.4 STA_VDBB.scala 326:29:@25006.4 STA_VDBB.scala 326:29:@25031.4 STA_VDBB.scala 326:29:@25798.4 STA_VDBB.scala 326:29:@25823.4 STA_VDBB.scala 326:29:@26590.4 STA_VDBB.scala 326:29:@26615.4 STA_VDBB.scala 326:29:@27382.4 STA_VDBB.scala 326:29:@27407.4]
  assign ff01_io_in_tag_2_6 = S8DP1_26_io_out_tag_6; // @[STA_VDBB.scala 109:23:@10242.4 STA_VDBB.scala 194:29:@13007.4 STA_VDBB.scala 194:29:@13032.4 STA_VDBB.scala 194:29:@13799.4 STA_VDBB.scala 194:29:@13824.4 STA_VDBB.scala 194:29:@14591.4 STA_VDBB.scala 194:29:@14616.4 STA_VDBB.scala 194:29:@15383.4 STA_VDBB.scala 194:29:@15408.4 STA_VDBB.scala 194:29:@16175.4 STA_VDBB.scala 194:29:@16200.4 STA_VDBB.scala 194:29:@16967.4 STA_VDBB.scala 194:29:@16992.4 STA_VDBB.scala 194:29:@17759.4 STA_VDBB.scala 194:29:@17784.4 STA_VDBB.scala 194:29:@18551.4 STA_VDBB.scala 194:29:@18576.4 STA_VDBB.scala 242:23:@19074.4 STA_VDBB.scala 326:29:@21839.4 STA_VDBB.scala 326:29:@21864.4 STA_VDBB.scala 326:29:@22631.4 STA_VDBB.scala 326:29:@22656.4 STA_VDBB.scala 326:29:@23423.4 STA_VDBB.scala 326:29:@23448.4 STA_VDBB.scala 326:29:@24215.4 STA_VDBB.scala 326:29:@24240.4 STA_VDBB.scala 326:29:@25007.4 STA_VDBB.scala 326:29:@25032.4 STA_VDBB.scala 326:29:@25799.4 STA_VDBB.scala 326:29:@25824.4 STA_VDBB.scala 326:29:@26591.4 STA_VDBB.scala 326:29:@26616.4 STA_VDBB.scala 326:29:@27383.4 STA_VDBB.scala 326:29:@27408.4]
  assign ff01_io_in_tag_2_7 = S8DP1_26_io_out_tag_7; // @[STA_VDBB.scala 109:23:@10243.4 STA_VDBB.scala 194:29:@13008.4 STA_VDBB.scala 194:29:@13033.4 STA_VDBB.scala 194:29:@13800.4 STA_VDBB.scala 194:29:@13825.4 STA_VDBB.scala 194:29:@14592.4 STA_VDBB.scala 194:29:@14617.4 STA_VDBB.scala 194:29:@15384.4 STA_VDBB.scala 194:29:@15409.4 STA_VDBB.scala 194:29:@16176.4 STA_VDBB.scala 194:29:@16201.4 STA_VDBB.scala 194:29:@16968.4 STA_VDBB.scala 194:29:@16993.4 STA_VDBB.scala 194:29:@17760.4 STA_VDBB.scala 194:29:@17785.4 STA_VDBB.scala 194:29:@18552.4 STA_VDBB.scala 194:29:@18577.4 STA_VDBB.scala 242:23:@19075.4 STA_VDBB.scala 326:29:@21840.4 STA_VDBB.scala 326:29:@21865.4 STA_VDBB.scala 326:29:@22632.4 STA_VDBB.scala 326:29:@22657.4 STA_VDBB.scala 326:29:@23424.4 STA_VDBB.scala 326:29:@23449.4 STA_VDBB.scala 326:29:@24216.4 STA_VDBB.scala 326:29:@24241.4 STA_VDBB.scala 326:29:@25008.4 STA_VDBB.scala 326:29:@25033.4 STA_VDBB.scala 326:29:@25800.4 STA_VDBB.scala 326:29:@25825.4 STA_VDBB.scala 326:29:@26592.4 STA_VDBB.scala 326:29:@26617.4 STA_VDBB.scala 326:29:@27384.4 STA_VDBB.scala 326:29:@27409.4]
  assign ff01_io_in_tag_3_0 = S8DP1_27_io_out_tag_0; // @[STA_VDBB.scala 109:23:@10260.4 STA_VDBB.scala 194:29:@13067.4 STA_VDBB.scala 194:29:@13092.4 STA_VDBB.scala 194:29:@13859.4 STA_VDBB.scala 194:29:@13884.4 STA_VDBB.scala 194:29:@14651.4 STA_VDBB.scala 194:29:@14676.4 STA_VDBB.scala 194:29:@15443.4 STA_VDBB.scala 194:29:@15468.4 STA_VDBB.scala 194:29:@16235.4 STA_VDBB.scala 194:29:@16260.4 STA_VDBB.scala 194:29:@17027.4 STA_VDBB.scala 194:29:@17052.4 STA_VDBB.scala 194:29:@17819.4 STA_VDBB.scala 194:29:@17844.4 STA_VDBB.scala 194:29:@18611.4 STA_VDBB.scala 194:29:@18636.4 STA_VDBB.scala 242:23:@19092.4 STA_VDBB.scala 326:29:@21899.4 STA_VDBB.scala 326:29:@21924.4 STA_VDBB.scala 326:29:@22691.4 STA_VDBB.scala 326:29:@22716.4 STA_VDBB.scala 326:29:@23483.4 STA_VDBB.scala 326:29:@23508.4 STA_VDBB.scala 326:29:@24275.4 STA_VDBB.scala 326:29:@24300.4 STA_VDBB.scala 326:29:@25067.4 STA_VDBB.scala 326:29:@25092.4 STA_VDBB.scala 326:29:@25859.4 STA_VDBB.scala 326:29:@25884.4 STA_VDBB.scala 326:29:@26651.4 STA_VDBB.scala 326:29:@26676.4 STA_VDBB.scala 326:29:@27443.4 STA_VDBB.scala 326:29:@27468.4]
  assign ff01_io_in_tag_3_1 = S8DP1_27_io_out_tag_1; // @[STA_VDBB.scala 109:23:@10261.4 STA_VDBB.scala 194:29:@13068.4 STA_VDBB.scala 194:29:@13093.4 STA_VDBB.scala 194:29:@13860.4 STA_VDBB.scala 194:29:@13885.4 STA_VDBB.scala 194:29:@14652.4 STA_VDBB.scala 194:29:@14677.4 STA_VDBB.scala 194:29:@15444.4 STA_VDBB.scala 194:29:@15469.4 STA_VDBB.scala 194:29:@16236.4 STA_VDBB.scala 194:29:@16261.4 STA_VDBB.scala 194:29:@17028.4 STA_VDBB.scala 194:29:@17053.4 STA_VDBB.scala 194:29:@17820.4 STA_VDBB.scala 194:29:@17845.4 STA_VDBB.scala 194:29:@18612.4 STA_VDBB.scala 194:29:@18637.4 STA_VDBB.scala 242:23:@19093.4 STA_VDBB.scala 326:29:@21900.4 STA_VDBB.scala 326:29:@21925.4 STA_VDBB.scala 326:29:@22692.4 STA_VDBB.scala 326:29:@22717.4 STA_VDBB.scala 326:29:@23484.4 STA_VDBB.scala 326:29:@23509.4 STA_VDBB.scala 326:29:@24276.4 STA_VDBB.scala 326:29:@24301.4 STA_VDBB.scala 326:29:@25068.4 STA_VDBB.scala 326:29:@25093.4 STA_VDBB.scala 326:29:@25860.4 STA_VDBB.scala 326:29:@25885.4 STA_VDBB.scala 326:29:@26652.4 STA_VDBB.scala 326:29:@26677.4 STA_VDBB.scala 326:29:@27444.4 STA_VDBB.scala 326:29:@27469.4]
  assign ff01_io_in_tag_3_2 = S8DP1_27_io_out_tag_2; // @[STA_VDBB.scala 109:23:@10262.4 STA_VDBB.scala 194:29:@13069.4 STA_VDBB.scala 194:29:@13094.4 STA_VDBB.scala 194:29:@13861.4 STA_VDBB.scala 194:29:@13886.4 STA_VDBB.scala 194:29:@14653.4 STA_VDBB.scala 194:29:@14678.4 STA_VDBB.scala 194:29:@15445.4 STA_VDBB.scala 194:29:@15470.4 STA_VDBB.scala 194:29:@16237.4 STA_VDBB.scala 194:29:@16262.4 STA_VDBB.scala 194:29:@17029.4 STA_VDBB.scala 194:29:@17054.4 STA_VDBB.scala 194:29:@17821.4 STA_VDBB.scala 194:29:@17846.4 STA_VDBB.scala 194:29:@18613.4 STA_VDBB.scala 194:29:@18638.4 STA_VDBB.scala 242:23:@19094.4 STA_VDBB.scala 326:29:@21901.4 STA_VDBB.scala 326:29:@21926.4 STA_VDBB.scala 326:29:@22693.4 STA_VDBB.scala 326:29:@22718.4 STA_VDBB.scala 326:29:@23485.4 STA_VDBB.scala 326:29:@23510.4 STA_VDBB.scala 326:29:@24277.4 STA_VDBB.scala 326:29:@24302.4 STA_VDBB.scala 326:29:@25069.4 STA_VDBB.scala 326:29:@25094.4 STA_VDBB.scala 326:29:@25861.4 STA_VDBB.scala 326:29:@25886.4 STA_VDBB.scala 326:29:@26653.4 STA_VDBB.scala 326:29:@26678.4 STA_VDBB.scala 326:29:@27445.4 STA_VDBB.scala 326:29:@27470.4]
  assign ff01_io_in_tag_3_3 = S8DP1_27_io_out_tag_3; // @[STA_VDBB.scala 109:23:@10263.4 STA_VDBB.scala 194:29:@13070.4 STA_VDBB.scala 194:29:@13095.4 STA_VDBB.scala 194:29:@13862.4 STA_VDBB.scala 194:29:@13887.4 STA_VDBB.scala 194:29:@14654.4 STA_VDBB.scala 194:29:@14679.4 STA_VDBB.scala 194:29:@15446.4 STA_VDBB.scala 194:29:@15471.4 STA_VDBB.scala 194:29:@16238.4 STA_VDBB.scala 194:29:@16263.4 STA_VDBB.scala 194:29:@17030.4 STA_VDBB.scala 194:29:@17055.4 STA_VDBB.scala 194:29:@17822.4 STA_VDBB.scala 194:29:@17847.4 STA_VDBB.scala 194:29:@18614.4 STA_VDBB.scala 194:29:@18639.4 STA_VDBB.scala 242:23:@19095.4 STA_VDBB.scala 326:29:@21902.4 STA_VDBB.scala 326:29:@21927.4 STA_VDBB.scala 326:29:@22694.4 STA_VDBB.scala 326:29:@22719.4 STA_VDBB.scala 326:29:@23486.4 STA_VDBB.scala 326:29:@23511.4 STA_VDBB.scala 326:29:@24278.4 STA_VDBB.scala 326:29:@24303.4 STA_VDBB.scala 326:29:@25070.4 STA_VDBB.scala 326:29:@25095.4 STA_VDBB.scala 326:29:@25862.4 STA_VDBB.scala 326:29:@25887.4 STA_VDBB.scala 326:29:@26654.4 STA_VDBB.scala 326:29:@26679.4 STA_VDBB.scala 326:29:@27446.4 STA_VDBB.scala 326:29:@27471.4]
  assign ff01_io_in_tag_3_4 = S8DP1_27_io_out_tag_4; // @[STA_VDBB.scala 109:23:@10264.4 STA_VDBB.scala 194:29:@13071.4 STA_VDBB.scala 194:29:@13096.4 STA_VDBB.scala 194:29:@13863.4 STA_VDBB.scala 194:29:@13888.4 STA_VDBB.scala 194:29:@14655.4 STA_VDBB.scala 194:29:@14680.4 STA_VDBB.scala 194:29:@15447.4 STA_VDBB.scala 194:29:@15472.4 STA_VDBB.scala 194:29:@16239.4 STA_VDBB.scala 194:29:@16264.4 STA_VDBB.scala 194:29:@17031.4 STA_VDBB.scala 194:29:@17056.4 STA_VDBB.scala 194:29:@17823.4 STA_VDBB.scala 194:29:@17848.4 STA_VDBB.scala 194:29:@18615.4 STA_VDBB.scala 194:29:@18640.4 STA_VDBB.scala 242:23:@19096.4 STA_VDBB.scala 326:29:@21903.4 STA_VDBB.scala 326:29:@21928.4 STA_VDBB.scala 326:29:@22695.4 STA_VDBB.scala 326:29:@22720.4 STA_VDBB.scala 326:29:@23487.4 STA_VDBB.scala 326:29:@23512.4 STA_VDBB.scala 326:29:@24279.4 STA_VDBB.scala 326:29:@24304.4 STA_VDBB.scala 326:29:@25071.4 STA_VDBB.scala 326:29:@25096.4 STA_VDBB.scala 326:29:@25863.4 STA_VDBB.scala 326:29:@25888.4 STA_VDBB.scala 326:29:@26655.4 STA_VDBB.scala 326:29:@26680.4 STA_VDBB.scala 326:29:@27447.4 STA_VDBB.scala 326:29:@27472.4]
  assign ff01_io_in_tag_3_5 = S8DP1_27_io_out_tag_5; // @[STA_VDBB.scala 109:23:@10265.4 STA_VDBB.scala 194:29:@13072.4 STA_VDBB.scala 194:29:@13097.4 STA_VDBB.scala 194:29:@13864.4 STA_VDBB.scala 194:29:@13889.4 STA_VDBB.scala 194:29:@14656.4 STA_VDBB.scala 194:29:@14681.4 STA_VDBB.scala 194:29:@15448.4 STA_VDBB.scala 194:29:@15473.4 STA_VDBB.scala 194:29:@16240.4 STA_VDBB.scala 194:29:@16265.4 STA_VDBB.scala 194:29:@17032.4 STA_VDBB.scala 194:29:@17057.4 STA_VDBB.scala 194:29:@17824.4 STA_VDBB.scala 194:29:@17849.4 STA_VDBB.scala 194:29:@18616.4 STA_VDBB.scala 194:29:@18641.4 STA_VDBB.scala 242:23:@19097.4 STA_VDBB.scala 326:29:@21904.4 STA_VDBB.scala 326:29:@21929.4 STA_VDBB.scala 326:29:@22696.4 STA_VDBB.scala 326:29:@22721.4 STA_VDBB.scala 326:29:@23488.4 STA_VDBB.scala 326:29:@23513.4 STA_VDBB.scala 326:29:@24280.4 STA_VDBB.scala 326:29:@24305.4 STA_VDBB.scala 326:29:@25072.4 STA_VDBB.scala 326:29:@25097.4 STA_VDBB.scala 326:29:@25864.4 STA_VDBB.scala 326:29:@25889.4 STA_VDBB.scala 326:29:@26656.4 STA_VDBB.scala 326:29:@26681.4 STA_VDBB.scala 326:29:@27448.4 STA_VDBB.scala 326:29:@27473.4]
  assign ff01_io_in_tag_3_6 = S8DP1_27_io_out_tag_6; // @[STA_VDBB.scala 109:23:@10266.4 STA_VDBB.scala 194:29:@13073.4 STA_VDBB.scala 194:29:@13098.4 STA_VDBB.scala 194:29:@13865.4 STA_VDBB.scala 194:29:@13890.4 STA_VDBB.scala 194:29:@14657.4 STA_VDBB.scala 194:29:@14682.4 STA_VDBB.scala 194:29:@15449.4 STA_VDBB.scala 194:29:@15474.4 STA_VDBB.scala 194:29:@16241.4 STA_VDBB.scala 194:29:@16266.4 STA_VDBB.scala 194:29:@17033.4 STA_VDBB.scala 194:29:@17058.4 STA_VDBB.scala 194:29:@17825.4 STA_VDBB.scala 194:29:@17850.4 STA_VDBB.scala 194:29:@18617.4 STA_VDBB.scala 194:29:@18642.4 STA_VDBB.scala 242:23:@19098.4 STA_VDBB.scala 326:29:@21905.4 STA_VDBB.scala 326:29:@21930.4 STA_VDBB.scala 326:29:@22697.4 STA_VDBB.scala 326:29:@22722.4 STA_VDBB.scala 326:29:@23489.4 STA_VDBB.scala 326:29:@23514.4 STA_VDBB.scala 326:29:@24281.4 STA_VDBB.scala 326:29:@24306.4 STA_VDBB.scala 326:29:@25073.4 STA_VDBB.scala 326:29:@25098.4 STA_VDBB.scala 326:29:@25865.4 STA_VDBB.scala 326:29:@25890.4 STA_VDBB.scala 326:29:@26657.4 STA_VDBB.scala 326:29:@26682.4 STA_VDBB.scala 326:29:@27449.4 STA_VDBB.scala 326:29:@27474.4]
  assign ff01_io_in_tag_3_7 = S8DP1_27_io_out_tag_7; // @[STA_VDBB.scala 109:23:@10267.4 STA_VDBB.scala 194:29:@13074.4 STA_VDBB.scala 194:29:@13099.4 STA_VDBB.scala 194:29:@13866.4 STA_VDBB.scala 194:29:@13891.4 STA_VDBB.scala 194:29:@14658.4 STA_VDBB.scala 194:29:@14683.4 STA_VDBB.scala 194:29:@15450.4 STA_VDBB.scala 194:29:@15475.4 STA_VDBB.scala 194:29:@16242.4 STA_VDBB.scala 194:29:@16267.4 STA_VDBB.scala 194:29:@17034.4 STA_VDBB.scala 194:29:@17059.4 STA_VDBB.scala 194:29:@17826.4 STA_VDBB.scala 194:29:@17851.4 STA_VDBB.scala 194:29:@18618.4 STA_VDBB.scala 194:29:@18643.4 STA_VDBB.scala 242:23:@19099.4 STA_VDBB.scala 326:29:@21906.4 STA_VDBB.scala 326:29:@21931.4 STA_VDBB.scala 326:29:@22698.4 STA_VDBB.scala 326:29:@22723.4 STA_VDBB.scala 326:29:@23490.4 STA_VDBB.scala 326:29:@23515.4 STA_VDBB.scala 326:29:@24282.4 STA_VDBB.scala 326:29:@24307.4 STA_VDBB.scala 326:29:@25074.4 STA_VDBB.scala 326:29:@25099.4 STA_VDBB.scala 326:29:@25866.4 STA_VDBB.scala 326:29:@25891.4 STA_VDBB.scala 326:29:@26658.4 STA_VDBB.scala 326:29:@26683.4 STA_VDBB.scala 326:29:@27450.4 STA_VDBB.scala 326:29:@27475.4]
  assign ff10_clock = clock; // @[:@9802.4]
  assign ff10_reset = reset; // @[:@9803.4]
  assign ff10_io_in_data_0_0 = io_in_B_4_8; // @[STA_VDBB.scala 154:29:@12385.4 STA_VDBB.scala 286:29:@21217.4]
  assign ff10_io_in_data_0_1 = io_in_B_4_9; // @[STA_VDBB.scala 154:29:@12397.4 STA_VDBB.scala 286:29:@21229.4]
  assign ff10_io_in_data_0_2 = io_in_B_4_10; // @[STA_VDBB.scala 154:29:@12409.4 STA_VDBB.scala 286:29:@21241.4]
  assign ff10_io_in_data_0_3 = io_in_B_4_11; // @[STA_VDBB.scala 154:29:@12421.4 STA_VDBB.scala 286:29:@21253.4]
  assign ff10_io_in_data_0_4 = io_in_B_4_12; // @[STA_VDBB.scala 154:29:@12433.4 STA_VDBB.scala 286:29:@21265.4]
  assign ff10_io_in_data_0_5 = io_in_B_4_13; // @[STA_VDBB.scala 154:29:@12445.4 STA_VDBB.scala 286:29:@21277.4]
  assign ff10_io_in_data_0_6 = io_in_B_4_14; // @[STA_VDBB.scala 154:29:@12457.4 STA_VDBB.scala 286:29:@21289.4]
  assign ff10_io_in_data_0_7 = io_in_B_4_15; // @[STA_VDBB.scala 154:29:@12469.4 STA_VDBB.scala 286:29:@21301.4]
  assign ff10_io_in_data_1_0 = io_in_B_5_8; // @[STA_VDBB.scala 154:29:@12387.4 STA_VDBB.scala 286:29:@21219.4]
  assign ff10_io_in_data_1_1 = io_in_B_5_9; // @[STA_VDBB.scala 154:29:@12399.4 STA_VDBB.scala 286:29:@21231.4]
  assign ff10_io_in_data_1_2 = io_in_B_5_10; // @[STA_VDBB.scala 154:29:@12411.4 STA_VDBB.scala 286:29:@21243.4]
  assign ff10_io_in_data_1_3 = io_in_B_5_11; // @[STA_VDBB.scala 154:29:@12423.4 STA_VDBB.scala 286:29:@21255.4]
  assign ff10_io_in_data_1_4 = io_in_B_5_12; // @[STA_VDBB.scala 154:29:@12435.4 STA_VDBB.scala 286:29:@21267.4]
  assign ff10_io_in_data_1_5 = io_in_B_5_13; // @[STA_VDBB.scala 154:29:@12447.4 STA_VDBB.scala 286:29:@21279.4]
  assign ff10_io_in_data_1_6 = io_in_B_5_14; // @[STA_VDBB.scala 154:29:@12459.4 STA_VDBB.scala 286:29:@21291.4]
  assign ff10_io_in_data_1_7 = io_in_B_5_15; // @[STA_VDBB.scala 154:29:@12471.4 STA_VDBB.scala 286:29:@21303.4]
  assign ff10_io_in_data_2_0 = io_in_B_6_8; // @[STA_VDBB.scala 154:29:@12389.4 STA_VDBB.scala 286:29:@21221.4]
  assign ff10_io_in_data_2_1 = io_in_B_6_9; // @[STA_VDBB.scala 154:29:@12401.4 STA_VDBB.scala 286:29:@21233.4]
  assign ff10_io_in_data_2_2 = io_in_B_6_10; // @[STA_VDBB.scala 154:29:@12413.4 STA_VDBB.scala 286:29:@21245.4]
  assign ff10_io_in_data_2_3 = io_in_B_6_11; // @[STA_VDBB.scala 154:29:@12425.4 STA_VDBB.scala 286:29:@21257.4]
  assign ff10_io_in_data_2_4 = io_in_B_6_12; // @[STA_VDBB.scala 154:29:@12437.4 STA_VDBB.scala 286:29:@21269.4]
  assign ff10_io_in_data_2_5 = io_in_B_6_13; // @[STA_VDBB.scala 154:29:@12449.4 STA_VDBB.scala 286:29:@21281.4]
  assign ff10_io_in_data_2_6 = io_in_B_6_14; // @[STA_VDBB.scala 154:29:@12461.4 STA_VDBB.scala 286:29:@21293.4]
  assign ff10_io_in_data_2_7 = io_in_B_6_15; // @[STA_VDBB.scala 154:29:@12473.4 STA_VDBB.scala 286:29:@21305.4]
  assign ff10_io_in_data_3_0 = io_in_B_7_8; // @[STA_VDBB.scala 154:29:@12391.4 STA_VDBB.scala 286:29:@21223.4]
  assign ff10_io_in_data_3_1 = io_in_B_7_9; // @[STA_VDBB.scala 154:29:@12403.4 STA_VDBB.scala 286:29:@21235.4]
  assign ff10_io_in_data_3_2 = io_in_B_7_10; // @[STA_VDBB.scala 154:29:@12415.4 STA_VDBB.scala 286:29:@21247.4]
  assign ff10_io_in_data_3_3 = io_in_B_7_11; // @[STA_VDBB.scala 154:29:@12427.4 STA_VDBB.scala 286:29:@21259.4]
  assign ff10_io_in_data_3_4 = io_in_B_7_12; // @[STA_VDBB.scala 154:29:@12439.4 STA_VDBB.scala 286:29:@21271.4]
  assign ff10_io_in_data_3_5 = io_in_B_7_13; // @[STA_VDBB.scala 154:29:@12451.4 STA_VDBB.scala 286:29:@21283.4]
  assign ff10_io_in_data_3_6 = io_in_B_7_14; // @[STA_VDBB.scala 154:29:@12463.4 STA_VDBB.scala 286:29:@21295.4]
  assign ff10_io_in_data_3_7 = io_in_B_7_15; // @[STA_VDBB.scala 154:29:@12475.4 STA_VDBB.scala 286:29:@21307.4]
  assign ff10_io_in_tag_0_0 = tag_io_out_tag_0; // @[STA_VDBB.scala 162:23:@12492.4 STA_VDBB.scala 294:23:@21324.4]
  assign ff10_io_in_tag_0_1 = tag_io_out_tag_1; // @[STA_VDBB.scala 162:23:@12493.4 STA_VDBB.scala 294:23:@21325.4]
  assign ff10_io_in_tag_0_2 = tag_io_out_tag_2; // @[STA_VDBB.scala 162:23:@12494.4 STA_VDBB.scala 294:23:@21326.4]
  assign ff10_io_in_tag_0_3 = tag_io_out_tag_3; // @[STA_VDBB.scala 162:23:@12495.4 STA_VDBB.scala 294:23:@21327.4]
  assign ff10_io_in_tag_0_4 = tag_io_out_tag_4; // @[STA_VDBB.scala 162:23:@12496.4 STA_VDBB.scala 294:23:@21328.4]
  assign ff10_io_in_tag_0_5 = tag_io_out_tag_5; // @[STA_VDBB.scala 162:23:@12497.4 STA_VDBB.scala 294:23:@21329.4]
  assign ff10_io_in_tag_0_6 = tag_io_out_tag_6; // @[STA_VDBB.scala 162:23:@12498.4 STA_VDBB.scala 294:23:@21330.4]
  assign ff10_io_in_tag_0_7 = 1'h0; // @[STA_VDBB.scala 162:23:@12499.4 STA_VDBB.scala 294:23:@21331.4]
  assign ff10_io_in_tag_1_0 = tag_1_io_out_tag_0; // @[STA_VDBB.scala 162:23:@12516.4 STA_VDBB.scala 294:23:@21348.4]
  assign ff10_io_in_tag_1_1 = tag_1_io_out_tag_1; // @[STA_VDBB.scala 162:23:@12517.4 STA_VDBB.scala 294:23:@21349.4]
  assign ff10_io_in_tag_1_2 = tag_1_io_out_tag_2; // @[STA_VDBB.scala 162:23:@12518.4 STA_VDBB.scala 294:23:@21350.4]
  assign ff10_io_in_tag_1_3 = tag_1_io_out_tag_3; // @[STA_VDBB.scala 162:23:@12519.4 STA_VDBB.scala 294:23:@21351.4]
  assign ff10_io_in_tag_1_4 = tag_1_io_out_tag_4; // @[STA_VDBB.scala 162:23:@12520.4 STA_VDBB.scala 294:23:@21352.4]
  assign ff10_io_in_tag_1_5 = tag_1_io_out_tag_5; // @[STA_VDBB.scala 162:23:@12521.4 STA_VDBB.scala 294:23:@21353.4]
  assign ff10_io_in_tag_1_6 = tag_1_io_out_tag_6; // @[STA_VDBB.scala 162:23:@12522.4 STA_VDBB.scala 294:23:@21354.4]
  assign ff10_io_in_tag_1_7 = 1'h0; // @[STA_VDBB.scala 162:23:@12523.4 STA_VDBB.scala 294:23:@21355.4]
  assign ff10_io_in_tag_2_0 = tag_2_io_out_tag_0; // @[STA_VDBB.scala 162:23:@12540.4 STA_VDBB.scala 294:23:@21372.4]
  assign ff10_io_in_tag_2_1 = tag_2_io_out_tag_1; // @[STA_VDBB.scala 162:23:@12541.4 STA_VDBB.scala 294:23:@21373.4]
  assign ff10_io_in_tag_2_2 = tag_2_io_out_tag_2; // @[STA_VDBB.scala 162:23:@12542.4 STA_VDBB.scala 294:23:@21374.4]
  assign ff10_io_in_tag_2_3 = tag_2_io_out_tag_3; // @[STA_VDBB.scala 162:23:@12543.4 STA_VDBB.scala 294:23:@21375.4]
  assign ff10_io_in_tag_2_4 = tag_2_io_out_tag_4; // @[STA_VDBB.scala 162:23:@12544.4 STA_VDBB.scala 294:23:@21376.4]
  assign ff10_io_in_tag_2_5 = tag_2_io_out_tag_5; // @[STA_VDBB.scala 162:23:@12545.4 STA_VDBB.scala 294:23:@21377.4]
  assign ff10_io_in_tag_2_6 = tag_2_io_out_tag_6; // @[STA_VDBB.scala 162:23:@12546.4 STA_VDBB.scala 294:23:@21378.4]
  assign ff10_io_in_tag_2_7 = 1'h0; // @[STA_VDBB.scala 162:23:@12547.4 STA_VDBB.scala 294:23:@21379.4]
  assign ff10_io_in_tag_3_0 = tag_3_io_out_tag_0; // @[STA_VDBB.scala 162:23:@12564.4 STA_VDBB.scala 294:23:@21396.4]
  assign ff10_io_in_tag_3_1 = tag_3_io_out_tag_1; // @[STA_VDBB.scala 162:23:@12565.4 STA_VDBB.scala 294:23:@21397.4]
  assign ff10_io_in_tag_3_2 = tag_3_io_out_tag_2; // @[STA_VDBB.scala 162:23:@12566.4 STA_VDBB.scala 294:23:@21398.4]
  assign ff10_io_in_tag_3_3 = tag_3_io_out_tag_3; // @[STA_VDBB.scala 162:23:@12567.4 STA_VDBB.scala 294:23:@21399.4]
  assign ff10_io_in_tag_3_4 = tag_3_io_out_tag_4; // @[STA_VDBB.scala 162:23:@12568.4 STA_VDBB.scala 294:23:@21400.4]
  assign ff10_io_in_tag_3_5 = tag_3_io_out_tag_5; // @[STA_VDBB.scala 162:23:@12569.4 STA_VDBB.scala 294:23:@21401.4]
  assign ff10_io_in_tag_3_6 = tag_3_io_out_tag_6; // @[STA_VDBB.scala 162:23:@12570.4 STA_VDBB.scala 294:23:@21402.4]
  assign ff10_io_in_tag_3_7 = 1'h0; // @[STA_VDBB.scala 162:23:@12571.4 STA_VDBB.scala 294:23:@21403.4]
  assign ffa2_clock = clock; // @[:@9805.4]
  assign ffa2_reset = reset; // @[:@9806.4]
  assign ffa2_io_in_data_0_0 = io_in_A_2_8; // @[STA_VDBB.scala 143:29:@12380.4 STA_VDBB.scala 275:29:@21212.4]
  assign ffa2_io_in_data_0_1 = io_in_A_2_9; // @[STA_VDBB.scala 143:29:@12392.4 STA_VDBB.scala 275:29:@21224.4]
  assign ffa2_io_in_data_0_2 = io_in_A_2_10; // @[STA_VDBB.scala 143:29:@12404.4 STA_VDBB.scala 275:29:@21236.4]
  assign ffa2_io_in_data_0_3 = io_in_A_2_11; // @[STA_VDBB.scala 143:29:@12416.4 STA_VDBB.scala 275:29:@21248.4]
  assign ffa2_io_in_data_0_4 = io_in_A_2_12; // @[STA_VDBB.scala 143:29:@12428.4 STA_VDBB.scala 275:29:@21260.4]
  assign ffa2_io_in_data_0_5 = io_in_A_2_13; // @[STA_VDBB.scala 143:29:@12440.4 STA_VDBB.scala 275:29:@21272.4]
  assign ffa2_io_in_data_0_6 = io_in_A_2_14; // @[STA_VDBB.scala 143:29:@12452.4 STA_VDBB.scala 275:29:@21284.4]
  assign ffa2_io_in_data_0_7 = io_in_A_2_15; // @[STA_VDBB.scala 143:29:@12464.4 STA_VDBB.scala 275:29:@21296.4]
  assign ffa2_io_in_data_1_0 = io_in_A_3_8; // @[STA_VDBB.scala 143:29:@12382.4 STA_VDBB.scala 275:29:@21214.4]
  assign ffa2_io_in_data_1_1 = io_in_A_3_9; // @[STA_VDBB.scala 143:29:@12394.4 STA_VDBB.scala 275:29:@21226.4]
  assign ffa2_io_in_data_1_2 = io_in_A_3_10; // @[STA_VDBB.scala 143:29:@12406.4 STA_VDBB.scala 275:29:@21238.4]
  assign ffa2_io_in_data_1_3 = io_in_A_3_11; // @[STA_VDBB.scala 143:29:@12418.4 STA_VDBB.scala 275:29:@21250.4]
  assign ffa2_io_in_data_1_4 = io_in_A_3_12; // @[STA_VDBB.scala 143:29:@12430.4 STA_VDBB.scala 275:29:@21262.4]
  assign ffa2_io_in_data_1_5 = io_in_A_3_13; // @[STA_VDBB.scala 143:29:@12442.4 STA_VDBB.scala 275:29:@21274.4]
  assign ffa2_io_in_data_1_6 = io_in_A_3_14; // @[STA_VDBB.scala 143:29:@12454.4 STA_VDBB.scala 275:29:@21286.4]
  assign ffa2_io_in_data_1_7 = io_in_A_3_15; // @[STA_VDBB.scala 143:29:@12466.4 STA_VDBB.scala 275:29:@21298.4]
  assign ff11_clock = clock; // @[:@9808.4]
  assign ff11_reset = reset; // @[:@9809.4]
  assign ff11_io_in_data_0_0 = io_in_A_2_8; // @[STA_VDBB.scala 144:29:@12381.4 STA_VDBB.scala 276:29:@21213.4]
  assign ff11_io_in_data_0_1 = io_in_A_2_9; // @[STA_VDBB.scala 144:29:@12393.4 STA_VDBB.scala 276:29:@21225.4]
  assign ff11_io_in_data_0_2 = io_in_A_2_10; // @[STA_VDBB.scala 144:29:@12405.4 STA_VDBB.scala 276:29:@21237.4]
  assign ff11_io_in_data_0_3 = io_in_A_2_11; // @[STA_VDBB.scala 144:29:@12417.4 STA_VDBB.scala 276:29:@21249.4]
  assign ff11_io_in_data_0_4 = io_in_A_2_12; // @[STA_VDBB.scala 144:29:@12429.4 STA_VDBB.scala 276:29:@21261.4]
  assign ff11_io_in_data_0_5 = io_in_A_2_13; // @[STA_VDBB.scala 144:29:@12441.4 STA_VDBB.scala 276:29:@21273.4]
  assign ff11_io_in_data_0_6 = io_in_A_2_14; // @[STA_VDBB.scala 144:29:@12453.4 STA_VDBB.scala 276:29:@21285.4]
  assign ff11_io_in_data_0_7 = io_in_A_2_15; // @[STA_VDBB.scala 144:29:@12465.4 STA_VDBB.scala 276:29:@21297.4]
  assign ff11_io_in_data_1_0 = io_in_A_3_8; // @[STA_VDBB.scala 144:29:@12383.4 STA_VDBB.scala 276:29:@21215.4]
  assign ff11_io_in_data_1_1 = io_in_A_3_9; // @[STA_VDBB.scala 144:29:@12395.4 STA_VDBB.scala 276:29:@21227.4]
  assign ff11_io_in_data_1_2 = io_in_A_3_10; // @[STA_VDBB.scala 144:29:@12407.4 STA_VDBB.scala 276:29:@21239.4]
  assign ff11_io_in_data_1_3 = io_in_A_3_11; // @[STA_VDBB.scala 144:29:@12419.4 STA_VDBB.scala 276:29:@21251.4]
  assign ff11_io_in_data_1_4 = io_in_A_3_12; // @[STA_VDBB.scala 144:29:@12431.4 STA_VDBB.scala 276:29:@21263.4]
  assign ff11_io_in_data_1_5 = io_in_A_3_13; // @[STA_VDBB.scala 144:29:@12443.4 STA_VDBB.scala 276:29:@21275.4]
  assign ff11_io_in_data_1_6 = io_in_A_3_14; // @[STA_VDBB.scala 144:29:@12455.4 STA_VDBB.scala 276:29:@21287.4]
  assign ff11_io_in_data_1_7 = io_in_A_3_15; // @[STA_VDBB.scala 144:29:@12467.4 STA_VDBB.scala 276:29:@21299.4]
`ifdef RANDOMIZE_GARBAGE_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_INVALID_ASSIGN
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_REG_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE_MEM_INIT
`define RANDOMIZE
`endif
`ifdef RANDOMIZE
  integer initvar;
  initial begin
`ifndef verilator
  #0.002 begin end
`endif
`ifdef RANDOMIZE_REG_INIT
  _RAND_0 = {1{$random}};
  out_result_0_0 = _RAND_0[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_1 = {1{$random}};
  out_result_0_1 = _RAND_1[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_2 = {1{$random}};
  out_result_0_2 = _RAND_2[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_3 = {1{$random}};
  out_result_0_3 = _RAND_3[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_4 = {1{$random}};
  out_result_0_4 = _RAND_4[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_5 = {1{$random}};
  out_result_0_5 = _RAND_5[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_6 = {1{$random}};
  out_result_0_6 = _RAND_6[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_7 = {1{$random}};
  out_result_0_7 = _RAND_7[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_8 = {1{$random}};
  out_result_1_0 = _RAND_8[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_9 = {1{$random}};
  out_result_1_1 = _RAND_9[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_10 = {1{$random}};
  out_result_1_2 = _RAND_10[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_11 = {1{$random}};
  out_result_1_3 = _RAND_11[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_12 = {1{$random}};
  out_result_1_4 = _RAND_12[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_13 = {1{$random}};
  out_result_1_5 = _RAND_13[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_14 = {1{$random}};
  out_result_1_6 = _RAND_14[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_15 = {1{$random}};
  out_result_1_7 = _RAND_15[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_16 = {1{$random}};
  out_result_2_0 = _RAND_16[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_17 = {1{$random}};
  out_result_2_1 = _RAND_17[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_18 = {1{$random}};
  out_result_2_2 = _RAND_18[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_19 = {1{$random}};
  out_result_2_3 = _RAND_19[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_20 = {1{$random}};
  out_result_2_4 = _RAND_20[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_21 = {1{$random}};
  out_result_2_5 = _RAND_21[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_22 = {1{$random}};
  out_result_2_6 = _RAND_22[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_23 = {1{$random}};
  out_result_2_7 = _RAND_23[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_24 = {1{$random}};
  out_result_3_0 = _RAND_24[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_25 = {1{$random}};
  out_result_3_1 = _RAND_25[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_26 = {1{$random}};
  out_result_3_2 = _RAND_26[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_27 = {1{$random}};
  out_result_3_3 = _RAND_27[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_28 = {1{$random}};
  out_result_3_4 = _RAND_28[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_29 = {1{$random}};
  out_result_3_5 = _RAND_29[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_30 = {1{$random}};
  out_result_3_6 = _RAND_30[31:0];
`endif // RANDOMIZE_REG_INIT
`ifdef RANDOMIZE_REG_INIT
  _RAND_31 = {1{$random}};
  out_result_3_7 = _RAND_31[31:0];
`endif // RANDOMIZE_REG_INIT
  end
`endif // RANDOMIZE
  always @(posedge clock) begin
    if (reset) begin
      out_result_0_0 <= 32'sh0;
    end else begin
      out_result_0_0 <= S8DP1s_0_0_result;
    end
    if (reset) begin
      out_result_0_1 <= 32'sh0;
    end else begin
      out_result_0_1 <= S8DP1s_0_1_result;
    end
    if (reset) begin
      out_result_0_2 <= 32'sh0;
    end else begin
      out_result_0_2 <= S8DP1s_0_2_result;
    end
    if (reset) begin
      out_result_0_3 <= 32'sh0;
    end else begin
      out_result_0_3 <= S8DP1s_0_3_result;
    end
    if (reset) begin
      out_result_0_4 <= 32'sh0;
    end else begin
      out_result_0_4 <= S8DP1s_0_4_result;
    end
    if (reset) begin
      out_result_0_5 <= 32'sh0;
    end else begin
      out_result_0_5 <= S8DP1s_0_5_result;
    end
    if (reset) begin
      out_result_0_6 <= 32'sh0;
    end else begin
      out_result_0_6 <= S8DP1s_0_6_result;
    end
    if (reset) begin
      out_result_0_7 <= 32'sh0;
    end else begin
      out_result_0_7 <= S8DP1s_0_7_result;
    end
    if (reset) begin
      out_result_1_0 <= 32'sh0;
    end else begin
      out_result_1_0 <= S8DP1s_1_0_result;
    end
    if (reset) begin
      out_result_1_1 <= 32'sh0;
    end else begin
      out_result_1_1 <= S8DP1s_1_1_result;
    end
    if (reset) begin
      out_result_1_2 <= 32'sh0;
    end else begin
      out_result_1_2 <= S8DP1s_1_2_result;
    end
    if (reset) begin
      out_result_1_3 <= 32'sh0;
    end else begin
      out_result_1_3 <= S8DP1s_1_3_result;
    end
    if (reset) begin
      out_result_1_4 <= 32'sh0;
    end else begin
      out_result_1_4 <= S8DP1s_1_4_result;
    end
    if (reset) begin
      out_result_1_5 <= 32'sh0;
    end else begin
      out_result_1_5 <= S8DP1s_1_5_result;
    end
    if (reset) begin
      out_result_1_6 <= 32'sh0;
    end else begin
      out_result_1_6 <= S8DP1s_1_6_result;
    end
    if (reset) begin
      out_result_1_7 <= 32'sh0;
    end else begin
      out_result_1_7 <= S8DP1s_1_7_result;
    end
    if (reset) begin
      out_result_2_0 <= 32'sh0;
    end else begin
      out_result_2_0 <= S8DP1s_2_0_result;
    end
    if (reset) begin
      out_result_2_1 <= 32'sh0;
    end else begin
      out_result_2_1 <= S8DP1s_2_1_result;
    end
    if (reset) begin
      out_result_2_2 <= 32'sh0;
    end else begin
      out_result_2_2 <= S8DP1s_2_2_result;
    end
    if (reset) begin
      out_result_2_3 <= 32'sh0;
    end else begin
      out_result_2_3 <= S8DP1s_2_3_result;
    end
    if (reset) begin
      out_result_2_4 <= 32'sh0;
    end else begin
      out_result_2_4 <= S8DP1s_2_4_result;
    end
    if (reset) begin
      out_result_2_5 <= 32'sh0;
    end else begin
      out_result_2_5 <= S8DP1s_2_5_result;
    end
    if (reset) begin
      out_result_2_6 <= 32'sh0;
    end else begin
      out_result_2_6 <= S8DP1s_2_6_result;
    end
    if (reset) begin
      out_result_2_7 <= 32'sh0;
    end else begin
      out_result_2_7 <= S8DP1s_2_7_result;
    end
    if (reset) begin
      out_result_3_0 <= 32'sh0;
    end else begin
      out_result_3_0 <= S8DP1s_3_0_result;
    end
    if (reset) begin
      out_result_3_1 <= 32'sh0;
    end else begin
      out_result_3_1 <= S8DP1s_3_1_result;
    end
    if (reset) begin
      out_result_3_2 <= 32'sh0;
    end else begin
      out_result_3_2 <= S8DP1s_3_2_result;
    end
    if (reset) begin
      out_result_3_3 <= 32'sh0;
    end else begin
      out_result_3_3 <= S8DP1s_3_3_result;
    end
    if (reset) begin
      out_result_3_4 <= 32'sh0;
    end else begin
      out_result_3_4 <= S8DP1s_3_4_result;
    end
    if (reset) begin
      out_result_3_5 <= 32'sh0;
    end else begin
      out_result_3_5 <= S8DP1s_3_5_result;
    end
    if (reset) begin
      out_result_3_6 <= 32'sh0;
    end else begin
      out_result_3_6 <= S8DP1s_3_6_result;
    end
    if (reset) begin
      out_result_3_7 <= 32'sh0;
    end else begin
      out_result_3_7 <= S8DP1s_3_7_result;
    end
  end
endmodule
