module Mux8( // @[:@3.2]
  input         clock, // @[:@4.4]
  input         reset, // @[:@5.4]
  input  [31:0] io_int_in_0, // @[:@6.4]
  input  [31:0] io_int_in_1, // @[:@6.4]
  input  [31:0] io_int_in_2, // @[:@6.4]
  input  [31:0] io_int_in_3, // @[:@6.4]
  input  [31:0] io_int_in_4, // @[:@6.4]
  input  [31:0] io_int_in_5, // @[:@6.4]
  input  [31:0] io_int_in_6, // @[:@6.4]
  input  [31:0] io_int_in_7, // @[:@6.4]
  input         io_tag_0, // @[:@6.4]
  input         io_tag_1, // @[:@6.4]
  input         io_tag_2, // @[:@6.4]
  input         io_tag_3, // @[:@6.4]
  input         io_tag_4, // @[:@6.4]
  input         io_tag_5, // @[:@6.4]
  input         io_tag_6, // @[:@6.4]
  input         io_tag_7, // @[:@6.4]
  output [31:0] io_choice // @[:@6.4]
);
  wire [31:0] _T_62; // @[Mux.scala 19:72:@9.4]
  wire [31:0] _T_63; // @[Mux.scala 19:72:@10.4]
  wire [31:0] _T_66; // @[Mux.scala 19:72:@13.4]
  wire [31:0] _T_67; // @[Mux.scala 19:72:@14.4]
  wire [31:0] _T_70; // @[Mux.scala 19:72:@17.4]
  wire [31:0] _T_71; // @[Mux.scala 19:72:@18.4]
  wire [31:0] _T_74; // @[Mux.scala 19:72:@21.4]
  wire [31:0] _T_75; // @[Mux.scala 19:72:@22.4]
  wire [31:0] _T_78; // @[Mux.scala 19:72:@25.4]
  wire [31:0] _T_79; // @[Mux.scala 19:72:@26.4]
  wire [31:0] _T_82; // @[Mux.scala 19:72:@29.4]
  wire [31:0] _T_83; // @[Mux.scala 19:72:@30.4]
  wire [31:0] _T_86; // @[Mux.scala 19:72:@33.4]
  wire [31:0] _T_87; // @[Mux.scala 19:72:@34.4]
  wire [31:0] _T_90; // @[Mux.scala 19:72:@37.4]
  wire [31:0] _T_91; // @[Mux.scala 19:72:@38.4]
  wire [31:0] _T_93; // @[Mux.scala 19:72:@40.4]
  wire [31:0] _T_95; // @[Mux.scala 19:72:@41.4]
  wire [31:0] _T_97; // @[Mux.scala 19:72:@42.4]
  wire [31:0] _T_99; // @[Mux.scala 19:72:@43.4]
  wire [31:0] _T_101; // @[Mux.scala 19:72:@44.4]
  wire [31:0] _T_103; // @[Mux.scala 19:72:@45.4]
  wire [31:0] _T_105; // @[Mux.scala 19:72:@46.4]
  wire [31:0] _T_107; // @[Mux.scala 19:72:@47.4]
  wire [31:0] _T_108; // @[Mux.scala 19:72:@48.4]
  wire [31:0] _T_109; // @[Mux.scala 19:72:@49.4]
  wire [31:0] _T_110; // @[Mux.scala 19:72:@50.4]
  wire [31:0] _T_111; // @[Mux.scala 19:72:@51.4]
  wire [31:0] _T_112; // @[Mux.scala 19:72:@52.4]
  wire [31:0] _T_113; // @[Mux.scala 19:72:@53.4]
  wire [31:0] _T_114; // @[Mux.scala 19:72:@54.4]
  wire [31:0] _T_115; // @[Mux.scala 19:72:@55.4]
  wire [31:0] _T_116; // @[Mux.scala 19:72:@56.4]
  wire [31:0] _T_117; // @[Mux.scala 19:72:@57.4]
  wire [31:0] _T_118; // @[Mux.scala 19:72:@58.4]
  wire [31:0] _T_119; // @[Mux.scala 19:72:@59.4]
  wire [31:0] _T_120; // @[Mux.scala 19:72:@60.4]
  wire [31:0] _T_121; // @[Mux.scala 19:72:@61.4]
  wire [31:0] _T_124; // @[Mux.scala 19:72:@63.4]
  assign _T_62 = $unsigned(io_int_in_0); // @[Mux.scala 19:72:@9.4]
  assign _T_63 = $signed(_T_62); // @[Mux.scala 19:72:@10.4]
  assign _T_66 = $unsigned(io_int_in_1); // @[Mux.scala 19:72:@13.4]
  assign _T_67 = $signed(_T_66); // @[Mux.scala 19:72:@14.4]
  assign _T_70 = $unsigned(io_int_in_2); // @[Mux.scala 19:72:@17.4]
  assign _T_71 = $signed(_T_70); // @[Mux.scala 19:72:@18.4]
  assign _T_74 = $unsigned(io_int_in_3); // @[Mux.scala 19:72:@21.4]
  assign _T_75 = $signed(_T_74); // @[Mux.scala 19:72:@22.4]
  assign _T_78 = $unsigned(io_int_in_4); // @[Mux.scala 19:72:@25.4]
  assign _T_79 = $signed(_T_78); // @[Mux.scala 19:72:@26.4]
  assign _T_82 = $unsigned(io_int_in_5); // @[Mux.scala 19:72:@29.4]
  assign _T_83 = $signed(_T_82); // @[Mux.scala 19:72:@30.4]
  assign _T_86 = $unsigned(io_int_in_6); // @[Mux.scala 19:72:@33.4]
  assign _T_87 = $signed(_T_86); // @[Mux.scala 19:72:@34.4]
  assign _T_90 = $unsigned(io_int_in_7); // @[Mux.scala 19:72:@37.4]
  assign _T_91 = $signed(_T_90); // @[Mux.scala 19:72:@38.4]
  assign _T_93 = io_tag_0 ? $signed(_T_63) : $signed(32'sh0); // @[Mux.scala 19:72:@40.4]
  assign _T_95 = io_tag_1 ? $signed(_T_67) : $signed(32'sh0); // @[Mux.scala 19:72:@41.4]
  assign _T_97 = io_tag_2 ? $signed(_T_71) : $signed(32'sh0); // @[Mux.scala 19:72:@42.4]
  assign _T_99 = io_tag_3 ? $signed(_T_75) : $signed(32'sh0); // @[Mux.scala 19:72:@43.4]
  assign _T_101 = io_tag_4 ? $signed(_T_79) : $signed(32'sh0); // @[Mux.scala 19:72:@44.4]
  assign _T_103 = io_tag_5 ? $signed(_T_83) : $signed(32'sh0); // @[Mux.scala 19:72:@45.4]
  assign _T_105 = io_tag_6 ? $signed(_T_87) : $signed(32'sh0); // @[Mux.scala 19:72:@46.4]
  assign _T_107 = io_tag_7 ? $signed(_T_91) : $signed(32'sh0); // @[Mux.scala 19:72:@47.4]
  assign _T_108 = $signed(_T_93) | $signed(_T_95); // @[Mux.scala 19:72:@48.4]
  assign _T_109 = $signed(_T_108); // @[Mux.scala 19:72:@49.4]
  assign _T_110 = $signed(_T_109) | $signed(_T_97); // @[Mux.scala 19:72:@50.4]
  assign _T_111 = $signed(_T_110); // @[Mux.scala 19:72:@51.4]
  assign _T_112 = $signed(_T_111) | $signed(_T_99); // @[Mux.scala 19:72:@52.4]
  assign _T_113 = $signed(_T_112); // @[Mux.scala 19:72:@53.4]
  assign _T_114 = $signed(_T_113) | $signed(_T_101); // @[Mux.scala 19:72:@54.4]
  assign _T_115 = $signed(_T_114); // @[Mux.scala 19:72:@55.4]
  assign _T_116 = $signed(_T_115) | $signed(_T_103); // @[Mux.scala 19:72:@56.4]
  assign _T_117 = $signed(_T_116); // @[Mux.scala 19:72:@57.4]
  assign _T_118 = $signed(_T_117) | $signed(_T_105); // @[Mux.scala 19:72:@58.4]
  assign _T_119 = $signed(_T_118); // @[Mux.scala 19:72:@59.4]
  assign _T_120 = $signed(_T_119) | $signed(_T_107); // @[Mux.scala 19:72:@60.4]
  assign _T_121 = $signed(_T_120); // @[Mux.scala 19:72:@61.4]
  assign _T_124 = $unsigned(_T_121); // @[Mux.scala 19:72:@63.4]
  assign io_choice = $signed(_T_124); // @[Mux8.scala 40:13:@66.4]
endmodule
